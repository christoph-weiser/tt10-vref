VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_cw_vref
  CLASS BLOCK ;
  FOREIGN tt_um_cw_vref ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNADIFFAREA 4.640000 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNADIFFAREA 4.640000 ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 320.000000 ;
    ANTENNADIFFAREA 9.280000 ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNAGATEAREA 12.000000 ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[5]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 1439.971802 ;
    ANTENNADIFFAREA 616.904358 ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 150.062500 ;
    ANTENNADIFFAREA 1196.067749 ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 1439.971802 ;
    ANTENNADIFFAREA 616.904358 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.600 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 3.600 5.000 5.200 220.760 ;
    END
  END VGND
  PIN VAPWR
    ANTENNAGATEAREA 2912.000000 ;
    ANTENNADIFFAREA 2005.394531 ;
    PORT
      LAYER met4 ;
        RECT 6.200 5.000 7.800 220.760 ;
    END
  END VAPWR
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  OBS
      LAYER nwell ;
        RECT 3.250 220.980 103.675 223.480 ;
        RECT 3.250 5.750 5.750 220.980 ;
        RECT 8.935 180.290 45.725 212.250 ;
        RECT 48.860 187.290 56.700 210.740 ;
      LAYER pwell ;
        RECT 9.140 168.330 52.250 178.810 ;
      LAYER nwell ;
        RECT 62.865 170.855 99.075 217.105 ;
        RECT 101.175 182.070 103.675 220.980 ;
        RECT 108.240 216.015 153.520 220.985 ;
        RECT 108.240 203.045 153.520 214.015 ;
      LAYER pwell ;
        RECT 108.440 184.690 153.320 201.100 ;
      LAYER nwell ;
        RECT 164.960 200.075 239.400 201.680 ;
      LAYER pwell ;
        RECT 165.155 198.875 166.525 199.685 ;
        RECT 167.020 199.555 168.365 199.785 ;
        RECT 166.535 198.875 168.365 199.555 ;
        RECT 168.835 199.555 170.180 199.785 ;
        RECT 168.835 198.875 170.665 199.555 ;
        RECT 170.675 198.875 176.185 199.685 ;
        RECT 176.195 198.875 178.025 199.685 ;
        RECT 178.045 198.960 178.475 199.745 ;
        RECT 178.980 199.555 180.325 199.785 ;
        RECT 178.495 198.875 180.325 199.555 ;
        RECT 180.335 198.875 185.845 199.685 ;
        RECT 185.855 198.875 187.685 199.685 ;
        RECT 188.155 199.555 189.500 199.785 ;
        RECT 188.155 198.875 189.985 199.555 ;
        RECT 190.925 198.960 191.355 199.745 ;
        RECT 191.375 198.875 196.885 199.685 ;
        RECT 198.300 199.555 199.645 199.785 ;
        RECT 197.815 198.875 199.645 199.555 ;
        RECT 199.655 198.875 203.325 199.685 ;
        RECT 203.805 198.960 204.235 199.745 ;
        RECT 204.255 198.875 207.005 199.685 ;
        RECT 207.475 199.555 208.820 199.785 ;
        RECT 207.475 198.875 209.305 199.555 ;
        RECT 209.315 198.875 214.825 199.685 ;
        RECT 214.835 198.875 216.665 199.685 ;
        RECT 216.685 198.960 217.115 199.745 ;
        RECT 217.620 199.555 218.965 199.785 ;
        RECT 217.135 198.875 218.965 199.555 ;
        RECT 218.975 198.875 224.485 199.685 ;
        RECT 224.495 198.875 226.325 199.685 ;
        RECT 227.280 199.555 228.625 199.785 ;
        RECT 226.795 198.875 228.625 199.555 ;
        RECT 229.565 198.960 229.995 199.745 ;
        RECT 230.015 198.875 235.525 199.685 ;
        RECT 236.480 199.555 237.825 199.785 ;
        RECT 235.995 198.875 237.825 199.555 ;
        RECT 237.835 198.875 239.205 199.685 ;
        RECT 165.295 198.665 165.465 198.875 ;
        RECT 166.675 198.665 166.845 198.875 ;
        RECT 168.510 198.715 168.630 198.825 ;
        RECT 170.355 198.685 170.525 198.875 ;
        RECT 170.815 198.685 170.985 198.875 ;
        RECT 172.195 198.665 172.365 198.855 ;
        RECT 176.335 198.685 176.505 198.875 ;
        RECT 177.715 198.665 177.885 198.855 ;
        RECT 178.635 198.685 178.805 198.875 ;
        RECT 180.475 198.685 180.645 198.875 ;
        RECT 183.235 198.665 183.405 198.855 ;
        RECT 185.995 198.685 186.165 198.875 ;
        RECT 187.830 198.715 187.950 198.825 ;
        RECT 188.755 198.665 188.925 198.855 ;
        RECT 189.675 198.685 189.845 198.875 ;
        RECT 190.145 198.720 190.305 198.830 ;
        RECT 190.590 198.715 190.710 198.825 ;
        RECT 191.515 198.665 191.685 198.875 ;
        RECT 197.035 198.665 197.205 198.855 ;
        RECT 197.955 198.685 198.125 198.875 ;
        RECT 199.795 198.685 199.965 198.875 ;
        RECT 202.555 198.665 202.725 198.855 ;
        RECT 203.470 198.715 203.590 198.825 ;
        RECT 204.395 198.685 204.565 198.875 ;
        RECT 207.150 198.715 207.270 198.825 ;
        RECT 208.075 198.665 208.245 198.855 ;
        RECT 208.995 198.685 209.165 198.875 ;
        RECT 209.455 198.685 209.625 198.875 ;
        RECT 213.595 198.665 213.765 198.855 ;
        RECT 214.975 198.685 215.145 198.875 ;
        RECT 216.350 198.715 216.470 198.825 ;
        RECT 217.275 198.665 217.445 198.875 ;
        RECT 219.115 198.685 219.285 198.875 ;
        RECT 222.795 198.665 222.965 198.855 ;
        RECT 224.635 198.685 224.805 198.875 ;
        RECT 226.470 198.715 226.590 198.825 ;
        RECT 226.935 198.685 227.105 198.875 ;
        RECT 228.315 198.665 228.485 198.855 ;
        RECT 228.785 198.720 228.945 198.830 ;
        RECT 230.155 198.685 230.325 198.875 ;
        RECT 233.835 198.665 234.005 198.855 ;
        RECT 235.670 198.715 235.790 198.825 ;
        RECT 236.135 198.685 236.305 198.875 ;
        RECT 237.510 198.715 237.630 198.825 ;
        RECT 238.895 198.665 239.065 198.875 ;
        RECT 165.155 197.855 166.525 198.665 ;
        RECT 166.535 197.855 172.045 198.665 ;
        RECT 172.055 197.855 177.565 198.665 ;
        RECT 177.575 197.855 183.085 198.665 ;
        RECT 183.095 197.855 188.605 198.665 ;
        RECT 188.615 197.855 190.445 198.665 ;
        RECT 190.925 197.795 191.355 198.580 ;
        RECT 191.375 197.855 196.885 198.665 ;
        RECT 196.895 197.855 202.405 198.665 ;
        RECT 202.415 197.855 207.925 198.665 ;
        RECT 207.935 197.855 213.445 198.665 ;
        RECT 213.455 197.855 216.205 198.665 ;
        RECT 216.685 197.795 217.115 198.580 ;
        RECT 217.135 197.855 222.645 198.665 ;
        RECT 222.655 197.855 228.165 198.665 ;
        RECT 228.175 197.855 233.685 198.665 ;
        RECT 233.695 197.855 237.365 198.665 ;
        RECT 237.835 197.855 239.205 198.665 ;
      LAYER nwell ;
        RECT 164.960 194.635 239.400 197.465 ;
      LAYER pwell ;
        RECT 165.155 193.435 166.525 194.245 ;
        RECT 166.535 193.435 172.045 194.245 ;
        RECT 172.055 193.435 177.565 194.245 ;
        RECT 178.045 193.520 178.475 194.305 ;
        RECT 178.495 193.435 184.005 194.245 ;
        RECT 184.015 193.435 189.525 194.245 ;
        RECT 189.535 193.435 195.045 194.245 ;
        RECT 195.055 193.435 200.565 194.245 ;
        RECT 200.575 193.435 203.325 194.245 ;
        RECT 203.805 193.520 204.235 194.305 ;
        RECT 204.255 193.435 209.765 194.245 ;
        RECT 209.775 193.435 215.285 194.245 ;
        RECT 215.295 193.435 220.805 194.245 ;
        RECT 220.815 193.435 226.325 194.245 ;
        RECT 226.335 193.435 229.085 194.245 ;
        RECT 229.565 193.520 229.995 194.305 ;
        RECT 230.015 193.435 235.525 194.245 ;
        RECT 235.535 193.435 237.365 194.245 ;
        RECT 237.835 193.435 239.205 194.245 ;
        RECT 165.295 193.225 165.465 193.435 ;
        RECT 166.675 193.225 166.845 193.435 ;
        RECT 172.195 193.245 172.365 193.435 ;
        RECT 174.035 193.225 174.205 193.415 ;
        RECT 174.495 193.225 174.665 193.415 ;
        RECT 177.255 193.225 177.425 193.415 ;
        RECT 177.715 193.385 177.885 193.415 ;
        RECT 177.710 193.275 177.885 193.385 ;
        RECT 177.715 193.225 177.885 193.275 ;
        RECT 178.635 193.245 178.805 193.435 ;
        RECT 184.155 193.415 184.325 193.435 ;
        RECT 180.475 193.225 180.645 193.415 ;
        RECT 182.315 193.225 182.485 193.415 ;
        RECT 183.690 193.275 183.810 193.385 ;
        RECT 184.155 193.245 184.330 193.415 ;
        RECT 184.160 193.225 184.330 193.245 ;
        RECT 187.835 193.225 188.005 193.415 ;
        RECT 189.675 193.245 189.845 193.435 ;
        RECT 190.590 193.275 190.710 193.385 ;
        RECT 191.515 193.225 191.685 193.415 ;
        RECT 194.275 193.225 194.445 193.415 ;
        RECT 195.195 193.245 195.365 193.435 ;
        RECT 196.110 193.275 196.230 193.385 ;
        RECT 197.495 193.225 197.665 193.415 ;
        RECT 197.955 193.225 198.125 193.415 ;
        RECT 200.715 193.225 200.885 193.435 ;
        RECT 203.470 193.275 203.590 193.385 ;
        RECT 204.395 193.245 204.565 193.435 ;
        RECT 206.235 193.225 206.405 193.415 ;
        RECT 209.915 193.245 210.085 193.435 ;
        RECT 211.755 193.225 211.925 193.415 ;
        RECT 215.435 193.225 215.605 193.435 ;
        RECT 217.275 193.225 217.445 193.415 ;
        RECT 220.955 193.245 221.125 193.435 ;
        RECT 222.795 193.225 222.965 193.415 ;
        RECT 226.475 193.245 226.645 193.435 ;
        RECT 228.315 193.225 228.485 193.415 ;
        RECT 229.230 193.275 229.350 193.385 ;
        RECT 230.155 193.245 230.325 193.435 ;
        RECT 233.835 193.225 234.005 193.415 ;
        RECT 235.675 193.245 235.845 193.435 ;
        RECT 237.510 193.275 237.630 193.385 ;
        RECT 238.895 193.225 239.065 193.435 ;
        RECT 165.155 192.415 166.525 193.225 ;
        RECT 166.535 192.415 172.045 193.225 ;
        RECT 172.975 192.445 174.345 193.225 ;
        RECT 174.355 192.445 175.725 193.225 ;
        RECT 175.735 192.545 177.565 193.225 ;
        RECT 177.575 192.315 180.325 193.225 ;
        RECT 180.335 192.545 182.165 193.225 ;
        RECT 180.820 192.315 182.165 192.545 ;
        RECT 182.175 192.445 183.545 193.225 ;
        RECT 184.015 192.315 187.670 193.225 ;
        RECT 187.695 192.415 190.445 193.225 ;
        RECT 190.925 192.355 191.355 193.140 ;
        RECT 191.375 192.315 194.125 193.225 ;
        RECT 194.135 192.415 195.965 193.225 ;
        RECT 196.445 192.315 197.795 193.225 ;
        RECT 197.815 192.315 200.565 193.225 ;
        RECT 200.575 192.415 206.085 193.225 ;
        RECT 206.095 192.415 211.605 193.225 ;
        RECT 211.615 192.415 215.285 193.225 ;
        RECT 215.295 192.415 216.665 193.225 ;
        RECT 216.685 192.355 217.115 193.140 ;
        RECT 217.135 192.415 222.645 193.225 ;
        RECT 222.655 192.415 228.165 193.225 ;
        RECT 228.175 192.415 233.685 193.225 ;
        RECT 233.695 192.415 237.365 193.225 ;
        RECT 237.835 192.415 239.205 193.225 ;
      LAYER nwell ;
        RECT 164.960 189.195 239.400 192.025 ;
      LAYER pwell ;
        RECT 165.155 187.995 166.525 188.805 ;
        RECT 166.535 187.995 167.905 188.775 ;
        RECT 167.915 187.995 169.745 188.805 ;
        RECT 169.755 187.995 171.125 188.775 ;
        RECT 171.135 187.995 173.885 188.905 ;
        RECT 174.035 187.995 177.485 188.905 ;
        RECT 178.045 188.080 178.475 188.865 ;
        RECT 178.635 187.995 182.085 188.905 ;
        RECT 182.635 188.225 184.470 188.905 ;
        RECT 182.780 187.995 184.470 188.225 ;
        RECT 184.935 187.995 186.305 188.775 ;
        RECT 186.315 188.225 188.150 188.905 ;
        RECT 186.460 187.995 188.150 188.225 ;
        RECT 189.535 187.995 193.190 188.905 ;
        RECT 193.215 187.995 195.965 188.805 ;
        RECT 196.435 188.225 198.270 188.905 ;
        RECT 196.580 187.995 198.270 188.225 ;
        RECT 198.735 187.995 202.405 188.805 ;
        RECT 202.415 187.995 203.785 188.805 ;
        RECT 203.805 188.080 204.235 188.865 ;
        RECT 204.255 187.995 209.765 188.805 ;
        RECT 209.775 187.995 215.285 188.805 ;
        RECT 216.215 187.995 218.965 188.905 ;
        RECT 218.975 187.995 224.485 188.805 ;
        RECT 224.495 187.995 226.325 188.805 ;
        RECT 226.335 187.995 229.085 188.905 ;
        RECT 229.565 188.080 229.995 188.865 ;
        RECT 230.015 187.995 231.385 188.775 ;
        RECT 231.395 187.995 232.765 188.775 ;
        RECT 232.775 187.995 234.145 188.775 ;
        RECT 234.155 187.995 237.825 188.805 ;
        RECT 237.835 187.995 239.205 188.805 ;
        RECT 165.295 187.785 165.465 187.995 ;
        RECT 166.675 187.945 166.845 187.995 ;
        RECT 166.670 187.835 166.845 187.945 ;
        RECT 166.675 187.805 166.845 187.835 ;
        RECT 167.135 187.785 167.305 187.975 ;
        RECT 168.055 187.805 168.225 187.995 ;
        RECT 168.515 187.785 168.685 187.975 ;
        RECT 169.895 187.785 170.065 187.995 ;
        RECT 171.275 187.805 171.445 187.995 ;
        RECT 174.035 187.785 174.205 187.975 ;
        RECT 174.505 187.830 174.665 187.940 ;
        RECT 176.795 187.785 176.965 187.975 ;
        RECT 177.255 187.805 177.425 187.995 ;
        RECT 177.710 187.835 177.830 187.945 ;
        RECT 180.475 187.785 180.645 187.975 ;
        RECT 180.930 187.835 181.050 187.945 ;
        RECT 181.395 187.785 181.565 187.975 ;
        RECT 181.855 187.805 182.025 187.995 ;
        RECT 182.780 187.975 182.950 187.995 ;
        RECT 182.310 187.835 182.430 187.945 ;
        RECT 182.775 187.805 182.950 187.975 ;
        RECT 182.775 187.785 182.945 187.805 ;
        RECT 185.075 187.785 185.245 187.975 ;
        RECT 185.535 187.785 185.705 187.975 ;
        RECT 185.995 187.805 186.165 187.995 ;
        RECT 186.460 187.805 186.630 187.995 ;
        RECT 187.835 187.785 188.005 187.975 ;
        RECT 188.765 187.840 188.925 187.950 ;
        RECT 189.215 187.785 189.385 187.975 ;
        RECT 189.680 187.805 189.850 187.995 ;
        RECT 190.595 187.785 190.765 187.975 ;
        RECT 191.510 187.835 191.630 187.945 ;
        RECT 191.975 187.785 192.145 187.975 ;
        RECT 193.355 187.945 193.525 187.995 ;
        RECT 193.350 187.835 193.525 187.945 ;
        RECT 193.355 187.805 193.525 187.835 ;
        RECT 193.820 187.785 193.990 187.975 ;
        RECT 196.110 187.835 196.230 187.945 ;
        RECT 196.580 187.805 196.750 187.995 ;
        RECT 197.490 187.835 197.610 187.945 ;
        RECT 197.960 187.785 198.130 187.975 ;
        RECT 198.875 187.805 199.045 187.995 ;
        RECT 202.555 187.785 202.725 187.995 ;
        RECT 203.015 187.785 203.185 187.975 ;
        RECT 204.395 187.805 204.565 187.995 ;
        RECT 206.695 187.785 206.865 187.975 ;
        RECT 208.075 187.785 208.245 187.975 ;
        RECT 209.915 187.805 210.085 187.995 ;
        RECT 211.755 187.785 211.925 187.975 ;
        RECT 213.135 187.785 213.305 187.975 ;
        RECT 213.595 187.785 213.765 187.975 ;
        RECT 214.975 187.785 215.145 187.975 ;
        RECT 215.445 187.840 215.605 187.950 ;
        RECT 216.355 187.945 216.525 187.995 ;
        RECT 216.350 187.835 216.525 187.945 ;
        RECT 216.355 187.805 216.525 187.835 ;
        RECT 217.275 187.785 217.445 187.975 ;
        RECT 218.655 187.785 218.825 187.975 ;
        RECT 219.115 187.805 219.285 187.995 ;
        RECT 220.955 187.785 221.125 187.975 ;
        RECT 221.415 187.785 221.585 187.975 ;
        RECT 222.795 187.785 222.965 187.975 ;
        RECT 224.635 187.805 224.805 187.995 ;
        RECT 226.475 187.805 226.645 187.995 ;
        RECT 229.230 187.835 229.350 187.945 ;
        RECT 230.155 187.805 230.325 187.995 ;
        RECT 232.455 187.805 232.625 187.995 ;
        RECT 233.835 187.805 234.005 187.995 ;
        RECT 234.295 187.805 234.465 187.995 ;
        RECT 234.755 187.785 234.925 187.975 ;
        RECT 236.135 187.785 236.305 187.975 ;
        RECT 236.595 187.785 236.765 187.975 ;
        RECT 238.895 187.785 239.065 187.995 ;
        RECT 165.155 186.975 166.525 187.785 ;
        RECT 166.995 187.005 168.365 187.785 ;
        RECT 168.375 187.005 169.745 187.785 ;
        RECT 169.755 187.105 171.585 187.785 ;
        RECT 171.605 187.105 174.345 187.785 ;
        RECT 175.275 187.105 177.105 187.785 ;
        RECT 170.240 186.875 171.585 187.105 ;
        RECT 177.255 186.875 180.705 187.785 ;
        RECT 181.255 187.005 182.625 187.785 ;
        RECT 182.635 187.005 184.005 187.785 ;
        RECT 184.015 187.005 185.385 187.785 ;
        RECT 185.395 187.005 186.765 187.785 ;
        RECT 186.775 187.005 188.145 187.785 ;
        RECT 188.155 187.005 189.525 187.785 ;
        RECT 189.535 187.005 190.905 187.785 ;
        RECT 190.925 186.915 191.355 187.700 ;
        RECT 191.835 187.005 193.205 187.785 ;
        RECT 193.675 186.875 197.330 187.785 ;
        RECT 197.815 186.875 201.470 187.785 ;
        RECT 201.495 187.005 202.865 187.785 ;
        RECT 202.875 186.975 206.545 187.785 ;
        RECT 206.555 186.975 207.925 187.785 ;
        RECT 207.935 186.875 210.685 187.785 ;
        RECT 210.695 187.005 212.065 187.785 ;
        RECT 212.075 187.005 213.445 187.785 ;
        RECT 213.455 187.005 214.825 187.785 ;
        RECT 214.835 187.005 216.205 187.785 ;
        RECT 216.685 186.915 217.115 187.700 ;
        RECT 217.135 187.005 218.505 187.785 ;
        RECT 218.515 187.005 219.885 187.785 ;
        RECT 219.895 187.005 221.265 187.785 ;
        RECT 221.275 187.005 222.645 187.785 ;
        RECT 222.655 187.615 224.415 187.785 ;
        RECT 222.655 187.570 224.910 187.615 ;
        RECT 222.655 187.535 225.850 187.570 ;
        RECT 227.210 187.535 232.305 187.785 ;
        RECT 222.655 187.105 232.305 187.535 ;
        RECT 223.980 186.935 227.210 187.105 ;
        RECT 224.920 186.890 227.210 186.935 ;
        RECT 225.860 186.855 227.210 186.890 ;
        RECT 230.285 186.875 232.305 187.105 ;
        RECT 232.315 186.875 235.065 187.785 ;
        RECT 235.075 187.005 236.445 187.785 ;
        RECT 236.455 186.975 237.825 187.785 ;
        RECT 237.835 186.975 239.205 187.785 ;
        RECT 230.285 186.855 231.205 186.875 ;
      LAYER nwell ;
        RECT 164.960 183.755 239.400 186.585 ;
      LAYER pwell ;
        RECT 165.155 182.555 166.525 183.365 ;
        RECT 166.535 182.555 167.905 183.335 ;
        RECT 167.915 183.235 169.260 183.465 ;
        RECT 167.915 182.555 169.745 183.235 ;
        RECT 169.770 182.555 173.425 183.465 ;
        RECT 174.355 182.555 178.010 183.465 ;
        RECT 178.045 182.640 178.475 183.425 ;
        RECT 178.635 182.555 182.085 183.465 ;
        RECT 182.635 182.555 184.005 183.335 ;
        RECT 184.015 182.785 185.850 183.465 ;
        RECT 186.315 182.785 188.150 183.465 ;
        RECT 184.160 182.555 185.850 182.785 ;
        RECT 186.460 182.555 188.150 182.785 ;
        RECT 188.615 182.555 192.270 183.465 ;
        RECT 192.295 183.235 193.225 183.465 ;
        RECT 192.295 182.555 196.195 183.235 ;
        RECT 196.895 182.555 200.550 183.465 ;
        RECT 211.140 183.450 212.490 183.485 ;
        RECT 201.035 182.555 202.405 183.335 ;
        RECT 202.415 182.555 203.785 183.335 ;
        RECT 203.805 182.640 204.235 183.425 ;
        RECT 210.200 183.405 212.490 183.450 ;
        RECT 204.255 182.555 206.085 183.365 ;
        RECT 206.555 182.555 207.925 183.335 ;
        RECT 209.260 183.235 212.490 183.405 ;
        RECT 215.565 183.465 216.485 183.485 ;
        RECT 215.565 183.235 217.585 183.465 ;
        RECT 223.100 183.450 224.450 183.485 ;
        RECT 222.160 183.405 224.450 183.450 ;
        RECT 207.935 182.805 217.585 183.235 ;
        RECT 207.935 182.770 211.130 182.805 ;
        RECT 207.935 182.725 210.190 182.770 ;
        RECT 207.935 182.555 209.695 182.725 ;
        RECT 212.490 182.555 217.585 182.805 ;
        RECT 217.595 182.555 218.965 183.335 ;
        RECT 221.220 183.235 224.450 183.405 ;
        RECT 227.525 183.465 228.445 183.485 ;
        RECT 227.525 183.235 229.545 183.465 ;
        RECT 219.895 182.805 229.545 183.235 ;
        RECT 219.895 182.770 223.090 182.805 ;
        RECT 219.895 182.725 222.150 182.770 ;
        RECT 219.895 182.555 221.655 182.725 ;
        RECT 224.450 182.555 229.545 182.805 ;
        RECT 229.565 182.640 229.995 183.425 ;
        RECT 230.015 182.555 231.385 183.335 ;
        RECT 231.395 182.555 232.765 183.335 ;
        RECT 232.775 182.555 234.145 183.335 ;
        RECT 234.155 182.555 235.525 183.335 ;
        RECT 235.535 182.555 236.905 183.335 ;
        RECT 237.835 182.555 239.205 183.365 ;
        RECT 165.295 182.345 165.465 182.555 ;
        RECT 166.675 182.345 166.845 182.555 ;
        RECT 168.515 182.345 168.685 182.535 ;
        RECT 169.435 182.365 169.605 182.555 ;
        RECT 172.470 182.345 172.640 182.535 ;
        RECT 173.110 182.365 173.280 182.555 ;
        RECT 173.585 182.400 173.745 182.510 ;
        RECT 174.500 182.365 174.670 182.555 ;
        RECT 176.330 182.395 176.450 182.505 ;
        RECT 176.795 182.345 176.965 182.535 ;
        RECT 181.395 182.345 181.565 182.535 ;
        RECT 181.855 182.365 182.025 182.555 ;
        RECT 182.310 182.395 182.430 182.505 ;
        RECT 182.775 182.365 182.945 182.555 ;
        RECT 184.160 182.365 184.330 182.555 ;
        RECT 185.075 182.345 185.245 182.535 ;
        RECT 185.535 182.345 185.705 182.535 ;
        RECT 186.460 182.365 186.630 182.555 ;
        RECT 187.190 182.345 187.360 182.535 ;
        RECT 188.760 182.365 188.930 182.555 ;
        RECT 191.525 182.390 191.685 182.500 ;
        RECT 192.440 182.345 192.610 182.535 ;
        RECT 192.710 182.365 192.880 182.555 ;
        RECT 195.010 182.345 195.180 182.535 ;
        RECT 196.570 182.395 196.690 182.505 ;
        RECT 197.040 182.365 197.210 182.555 ;
        RECT 199.150 182.345 199.320 182.535 ;
        RECT 200.710 182.395 200.830 182.505 ;
        RECT 202.095 182.365 202.265 182.555 ;
        RECT 203.015 182.345 203.185 182.535 ;
        RECT 203.475 182.365 203.645 182.555 ;
        RECT 204.395 182.345 204.565 182.555 ;
        RECT 205.775 182.345 205.945 182.535 ;
        RECT 206.230 182.395 206.350 182.505 ;
        RECT 206.695 182.365 206.865 182.555 ;
        RECT 207.155 182.345 207.325 182.535 ;
        RECT 208.075 182.365 208.245 182.555 ;
        RECT 217.275 182.345 217.445 182.535 ;
        RECT 217.735 182.365 217.905 182.555 ;
        RECT 219.125 182.400 219.285 182.510 ;
        RECT 220.035 182.365 220.205 182.555 ;
        RECT 226.935 182.345 227.105 182.535 ;
        RECT 231.075 182.365 231.245 182.555 ;
        RECT 232.455 182.365 232.625 182.555 ;
        RECT 233.835 182.365 234.005 182.555 ;
        RECT 235.215 182.365 235.385 182.555 ;
        RECT 236.595 182.365 236.765 182.555 ;
        RECT 237.065 182.400 237.225 182.510 ;
        RECT 237.515 182.345 237.685 182.535 ;
        RECT 238.895 182.345 239.065 182.555 ;
      LAYER nwell ;
        RECT 101.175 179.570 156.750 182.070 ;
      LAYER pwell ;
        RECT 165.155 181.535 166.525 182.345 ;
        RECT 166.535 181.665 168.365 182.345 ;
        RECT 168.455 181.435 171.905 182.345 ;
        RECT 172.055 181.665 175.955 182.345 ;
        RECT 172.055 181.435 172.985 181.665 ;
        RECT 176.655 181.565 178.025 182.345 ;
        RECT 178.175 181.435 181.625 182.345 ;
        RECT 181.855 181.435 185.305 182.345 ;
        RECT 185.395 181.565 186.765 182.345 ;
        RECT 186.775 181.665 190.675 182.345 ;
        RECT 186.775 181.435 187.705 181.665 ;
        RECT 190.925 181.475 191.355 182.260 ;
        RECT 192.440 182.115 194.130 182.345 ;
        RECT 192.295 181.435 194.130 182.115 ;
        RECT 194.595 181.665 198.495 182.345 ;
        RECT 198.735 181.665 202.635 182.345 ;
        RECT 194.595 181.435 195.525 181.665 ;
        RECT 198.735 181.435 199.665 181.665 ;
        RECT 202.875 181.565 204.245 182.345 ;
        RECT 204.255 181.565 205.625 182.345 ;
        RECT 205.635 181.565 207.005 182.345 ;
        RECT 207.015 182.175 208.775 182.345 ;
        RECT 207.015 182.130 209.270 182.175 ;
        RECT 207.015 182.095 210.210 182.130 ;
        RECT 211.570 182.095 216.665 182.345 ;
        RECT 207.015 181.665 216.665 182.095 ;
        RECT 208.340 181.495 211.570 181.665 ;
        RECT 209.280 181.450 211.570 181.495 ;
        RECT 210.220 181.415 211.570 181.450 ;
        RECT 214.645 181.435 216.665 181.665 ;
        RECT 216.685 181.475 217.115 182.260 ;
        RECT 217.135 182.175 218.895 182.345 ;
        RECT 217.135 182.130 219.390 182.175 ;
        RECT 217.135 182.095 220.330 182.130 ;
        RECT 221.690 182.095 226.785 182.345 ;
        RECT 217.135 181.665 226.785 182.095 ;
        RECT 226.795 182.175 228.555 182.345 ;
        RECT 226.795 182.130 229.050 182.175 ;
        RECT 226.795 182.095 229.990 182.130 ;
        RECT 231.350 182.095 236.445 182.345 ;
        RECT 226.795 181.665 236.445 182.095 ;
        RECT 218.460 181.495 221.690 181.665 ;
        RECT 219.400 181.450 221.690 181.495 ;
        RECT 214.645 181.415 215.565 181.435 ;
        RECT 220.340 181.415 221.690 181.450 ;
        RECT 224.765 181.435 226.785 181.665 ;
        RECT 228.120 181.495 231.350 181.665 ;
        RECT 229.060 181.450 231.350 181.495 ;
        RECT 224.765 181.415 225.685 181.435 ;
        RECT 230.000 181.415 231.350 181.450 ;
        RECT 234.425 181.435 236.445 181.665 ;
        RECT 236.455 181.565 237.825 182.345 ;
        RECT 237.835 181.535 239.205 182.345 ;
        RECT 234.425 181.415 235.345 181.435 ;
        RECT 9.140 147.810 51.970 168.220 ;
      LAYER nwell ;
        RECT 63.050 164.975 97.990 167.475 ;
      LAYER pwell ;
        RECT 9.600 134.835 20.550 138.315 ;
        RECT 23.425 135.385 58.475 143.515 ;
      LAYER nwell ;
        RECT 63.050 135.035 65.550 164.975 ;
        RECT 69.300 160.385 91.740 161.225 ;
        RECT 69.300 139.625 70.140 160.385 ;
      LAYER pwell ;
        RECT 71.090 158.670 89.950 159.435 ;
        RECT 71.090 156.220 71.855 158.670 ;
        RECT 74.305 156.220 75.575 158.670 ;
        RECT 78.025 156.220 79.295 158.670 ;
        RECT 81.745 156.220 83.015 158.670 ;
        RECT 85.465 156.220 86.735 158.670 ;
        RECT 89.185 156.220 89.950 158.670 ;
        RECT 71.090 154.950 89.950 156.220 ;
        RECT 71.090 152.500 71.855 154.950 ;
        RECT 74.305 152.500 75.575 154.950 ;
        RECT 78.025 152.500 79.295 154.950 ;
        RECT 81.745 152.500 83.015 154.950 ;
        RECT 85.465 152.500 86.735 154.950 ;
        RECT 89.185 152.500 89.950 154.950 ;
        RECT 71.090 151.230 89.950 152.500 ;
        RECT 71.090 148.780 71.855 151.230 ;
        RECT 74.305 148.780 75.575 151.230 ;
        RECT 78.025 148.780 79.295 151.230 ;
        RECT 81.745 148.780 83.015 151.230 ;
        RECT 85.465 148.780 86.735 151.230 ;
        RECT 89.185 148.780 89.950 151.230 ;
        RECT 71.090 147.510 89.950 148.780 ;
        RECT 71.090 145.060 71.855 147.510 ;
        RECT 74.305 145.060 75.575 147.510 ;
        RECT 78.025 145.060 79.295 147.510 ;
        RECT 81.745 145.060 83.015 147.510 ;
        RECT 85.465 145.060 86.735 147.510 ;
        RECT 89.185 145.060 89.950 147.510 ;
        RECT 71.090 143.790 89.950 145.060 ;
        RECT 71.090 141.340 71.855 143.790 ;
        RECT 74.305 141.340 75.575 143.790 ;
        RECT 78.025 141.340 79.295 143.790 ;
        RECT 81.745 141.340 83.015 143.790 ;
        RECT 85.465 141.340 86.735 143.790 ;
        RECT 89.185 141.340 89.950 143.790 ;
        RECT 71.090 140.575 89.950 141.340 ;
      LAYER nwell ;
        RECT 90.900 139.625 91.740 160.385 ;
        RECT 69.300 138.785 91.740 139.625 ;
        RECT 95.490 135.035 97.990 164.975 ;
      LAYER pwell ;
        RECT 102.550 158.280 111.160 172.690 ;
        RECT 114.030 166.235 151.540 176.715 ;
      LAYER nwell ;
        RECT 102.350 141.345 111.360 156.335 ;
        RECT 115.985 139.690 149.475 158.060 ;
        RECT 63.050 132.535 97.990 135.035 ;
        RECT 138.080 129.720 145.960 134.690 ;
      LAYER pwell ;
        RECT 138.280 124.290 145.760 128.770 ;
      LAYER nwell ;
        RECT 10.025 41.635 128.935 124.285 ;
      LAYER pwell ;
        RECT 10.225 9.090 74.495 39.430 ;
        RECT 79.865 9.090 128.735 39.430 ;
      LAYER nwell ;
        RECT 135.120 13.460 149.570 109.050 ;
        RECT 154.250 5.750 156.750 179.570 ;
        RECT 164.960 178.315 239.400 181.145 ;
      LAYER pwell ;
        RECT 208.115 178.025 209.035 178.045 ;
        RECT 165.155 177.115 166.525 177.925 ;
        RECT 166.995 177.115 168.365 177.895 ;
        RECT 168.375 177.115 169.745 177.895 ;
        RECT 169.755 177.345 171.590 178.025 ;
        RECT 169.900 177.115 171.590 177.345 ;
        RECT 172.195 177.115 175.645 178.025 ;
        RECT 175.735 177.345 177.570 178.025 ;
        RECT 175.880 177.115 177.570 177.345 ;
        RECT 178.045 177.200 178.475 177.985 ;
        RECT 178.495 177.115 179.865 177.895 ;
        RECT 179.875 177.115 181.245 177.895 ;
        RECT 181.255 177.115 182.625 177.895 ;
        RECT 182.635 177.115 184.005 177.895 ;
        RECT 184.015 177.115 185.385 177.895 ;
        RECT 185.395 177.795 186.325 178.025 ;
        RECT 185.395 177.115 189.295 177.795 ;
        RECT 189.535 177.115 190.905 177.895 ;
        RECT 190.925 177.200 191.355 177.985 ;
        RECT 191.375 177.115 192.745 177.895 ;
        RECT 192.755 177.795 193.685 178.025 ;
        RECT 192.755 177.115 196.655 177.795 ;
        RECT 196.895 177.115 198.265 177.895 ;
        RECT 198.275 177.795 199.205 178.025 ;
        RECT 198.275 177.115 202.175 177.795 ;
        RECT 202.415 177.115 203.785 177.895 ;
        RECT 203.805 177.200 204.235 177.985 ;
        RECT 204.715 177.115 206.085 177.895 ;
        RECT 207.015 177.795 209.035 178.025 ;
        RECT 212.110 178.010 213.460 178.045 ;
        RECT 223.100 178.010 224.450 178.045 ;
        RECT 212.110 177.965 214.400 178.010 ;
        RECT 212.110 177.795 215.340 177.965 ;
        RECT 207.015 177.365 216.665 177.795 ;
        RECT 207.015 177.115 212.110 177.365 ;
        RECT 213.470 177.330 216.665 177.365 ;
        RECT 214.410 177.285 216.665 177.330 ;
        RECT 214.905 177.115 216.665 177.285 ;
        RECT 216.685 177.200 217.115 177.985 ;
        RECT 222.160 177.965 224.450 178.010 ;
        RECT 217.135 177.115 218.505 177.895 ;
        RECT 218.515 177.115 219.885 177.895 ;
        RECT 221.220 177.795 224.450 177.965 ;
        RECT 227.525 178.025 228.445 178.045 ;
        RECT 227.525 177.795 229.545 178.025 ;
        RECT 219.895 177.365 229.545 177.795 ;
        RECT 219.895 177.330 223.090 177.365 ;
        RECT 219.895 177.285 222.150 177.330 ;
        RECT 219.895 177.115 221.655 177.285 ;
        RECT 224.450 177.115 229.545 177.365 ;
        RECT 229.565 177.200 229.995 177.985 ;
        RECT 230.015 177.115 231.385 177.895 ;
        RECT 231.395 177.115 232.765 177.895 ;
        RECT 232.775 177.115 234.145 177.895 ;
        RECT 234.155 177.115 235.525 177.895 ;
        RECT 235.535 177.115 236.905 177.895 ;
        RECT 237.835 177.115 239.205 177.925 ;
        RECT 165.295 176.925 165.465 177.115 ;
        RECT 166.670 176.955 166.790 177.065 ;
        RECT 167.135 176.925 167.305 177.115 ;
        RECT 168.515 176.925 168.685 177.115 ;
        RECT 169.900 176.925 170.070 177.115 ;
        RECT 175.415 176.925 175.585 177.115 ;
        RECT 175.880 176.925 176.050 177.115 ;
        RECT 178.635 176.925 178.805 177.115 ;
        RECT 180.015 176.925 180.185 177.115 ;
        RECT 181.395 176.925 181.565 177.115 ;
        RECT 183.695 176.925 183.865 177.115 ;
        RECT 184.155 176.925 184.325 177.115 ;
        RECT 185.810 176.925 185.980 177.115 ;
        RECT 189.675 176.925 189.845 177.115 ;
        RECT 191.515 176.925 191.685 177.115 ;
        RECT 193.170 176.925 193.340 177.115 ;
        RECT 197.035 176.925 197.205 177.115 ;
        RECT 198.690 176.925 198.860 177.115 ;
        RECT 202.555 176.925 202.725 177.115 ;
        RECT 204.390 176.955 204.510 177.065 ;
        RECT 204.855 176.925 205.025 177.115 ;
        RECT 206.245 176.960 206.405 177.070 ;
        RECT 216.355 176.925 216.525 177.115 ;
        RECT 217.275 176.925 217.445 177.115 ;
        RECT 218.655 176.925 218.825 177.115 ;
        RECT 220.035 176.925 220.205 177.115 ;
        RECT 231.075 176.925 231.245 177.115 ;
        RECT 232.455 176.925 232.625 177.115 ;
        RECT 233.835 176.925 234.005 177.115 ;
        RECT 235.215 176.925 235.385 177.115 ;
        RECT 236.595 176.925 236.765 177.115 ;
        RECT 237.065 176.960 237.225 177.070 ;
        RECT 238.895 176.925 239.065 177.115 ;
        RECT 162.240 106.320 162.410 106.510 ;
        RECT 163.615 106.370 163.735 106.480 ;
        RECT 165.460 106.320 165.630 106.510 ;
        RECT 167.300 106.320 167.470 106.510 ;
        RECT 169.140 106.320 169.310 106.510 ;
        RECT 170.980 106.320 171.150 106.510 ;
        RECT 172.820 106.320 172.990 106.510 ;
        RECT 173.280 106.320 173.450 106.510 ;
        RECT 175.855 106.320 176.025 106.510 ;
        RECT 179.730 106.365 179.890 106.475 ;
        RECT 180.640 106.320 180.810 106.510 ;
        RECT 182.480 106.320 182.650 106.510 ;
        RECT 187.540 106.320 187.710 106.510 ;
        RECT 188.460 106.320 188.630 106.510 ;
        RECT 197.660 106.320 197.830 106.510 ;
        RECT 199.040 106.320 199.210 106.510 ;
        RECT 201.340 106.320 201.510 106.510 ;
        RECT 203.180 106.320 203.350 106.510 ;
        RECT 206.400 106.320 206.570 106.510 ;
        RECT 207.135 106.320 207.305 106.510 ;
        RECT 211.010 106.365 211.170 106.475 ;
        RECT 213.300 106.320 213.470 106.510 ;
        RECT 215.600 106.320 215.770 106.510 ;
        RECT 217.440 106.320 217.610 106.510 ;
        RECT 217.900 106.320 218.070 106.510 ;
        RECT 220.015 106.320 220.185 106.510 ;
        RECT 223.890 106.365 224.050 106.475 ;
        RECT 226.180 106.320 226.350 106.510 ;
        RECT 230.320 106.320 230.490 106.510 ;
        RECT 230.775 106.370 230.895 106.480 ;
        RECT 232.620 106.320 232.790 106.510 ;
        RECT 233.075 106.370 233.195 106.480 ;
        RECT 234.920 106.320 235.090 106.510 ;
        RECT 235.375 106.370 235.495 106.480 ;
        RECT 235.840 106.320 236.010 106.510 ;
        RECT 239.060 106.320 239.230 106.510 ;
        RECT 240.255 106.320 240.425 106.510 ;
        RECT 247.340 106.320 247.510 106.510 ;
        RECT 251.020 106.320 251.190 106.510 ;
        RECT 251.490 106.365 251.650 106.475 ;
        RECT 252.860 106.320 253.030 106.510 ;
        RECT 256.550 106.365 256.710 106.475 ;
        RECT 257.735 106.320 257.905 106.510 ;
        RECT 261.600 106.320 261.770 106.510 ;
        RECT 263.440 106.320 263.610 106.510 ;
        RECT 267.120 106.320 267.290 106.510 ;
        RECT 268.960 106.320 269.130 106.510 ;
        RECT 270.800 106.320 270.970 106.510 ;
        RECT 271.260 106.320 271.430 106.510 ;
        RECT 275.860 106.320 276.030 106.510 ;
        RECT 277.700 106.320 277.870 106.510 ;
        RECT 287.360 106.320 287.530 106.510 ;
        RECT 289.200 106.320 289.370 106.510 ;
        RECT 289.660 106.320 289.830 106.510 ;
        RECT 292.880 106.320 293.050 106.510 ;
        RECT 293.340 106.320 293.510 106.510 ;
        RECT 294.720 106.320 294.890 106.510 ;
        RECT 305.760 106.320 305.930 106.510 ;
        RECT 306.230 106.365 306.390 106.475 ;
        RECT 307.140 106.320 307.310 106.510 ;
        RECT 308.990 106.365 309.150 106.475 ;
        RECT 310.820 106.320 310.990 106.510 ;
        RECT 162.100 105.510 163.470 106.320 ;
        RECT 163.940 105.640 165.770 106.320 ;
        RECT 165.780 105.640 167.610 106.320 ;
        RECT 167.620 105.640 169.450 106.320 ;
        RECT 169.460 105.640 171.290 106.320 ;
        RECT 171.300 105.640 173.130 106.320 ;
        RECT 173.140 105.640 174.970 106.320 ;
        RECT 163.940 105.410 165.285 105.640 ;
        RECT 165.780 105.410 167.125 105.640 ;
        RECT 167.620 105.410 168.965 105.640 ;
        RECT 169.460 105.410 170.805 105.640 ;
        RECT 171.300 105.410 172.645 105.640 ;
        RECT 173.625 105.410 174.970 105.640 ;
        RECT 174.990 105.450 175.420 106.235 ;
        RECT 175.440 105.640 179.340 106.320 ;
        RECT 180.500 105.640 182.330 106.320 ;
        RECT 182.340 105.640 184.170 106.320 ;
        RECT 175.440 105.410 176.370 105.640 ;
        RECT 180.985 105.410 182.330 105.640 ;
        RECT 182.825 105.410 184.170 105.640 ;
        RECT 184.275 105.640 187.740 106.320 ;
        RECT 184.275 105.410 185.195 105.640 ;
        RECT 187.870 105.450 188.300 106.235 ;
        RECT 188.320 105.640 197.510 106.320 ;
        RECT 192.830 105.420 193.760 105.640 ;
        RECT 196.590 105.410 197.510 105.640 ;
        RECT 197.520 105.510 198.890 106.320 ;
        RECT 198.900 105.640 200.730 106.320 ;
        RECT 199.385 105.410 200.730 105.640 ;
        RECT 200.750 105.450 201.180 106.235 ;
        RECT 201.200 105.640 203.030 106.320 ;
        RECT 203.040 105.640 204.870 106.320 ;
        RECT 201.685 105.410 203.030 105.640 ;
        RECT 203.525 105.410 204.870 105.640 ;
        RECT 204.880 105.640 206.710 106.320 ;
        RECT 206.720 105.640 210.620 106.320 ;
        RECT 211.780 105.640 213.610 106.320 ;
        RECT 204.880 105.410 206.225 105.640 ;
        RECT 206.720 105.410 207.650 105.640 ;
        RECT 211.780 105.410 213.125 105.640 ;
        RECT 213.630 105.450 214.060 106.235 ;
        RECT 214.080 105.640 215.910 106.320 ;
        RECT 215.920 105.640 217.750 106.320 ;
        RECT 217.760 105.640 219.590 106.320 ;
        RECT 214.080 105.410 215.425 105.640 ;
        RECT 215.920 105.410 217.265 105.640 ;
        RECT 218.245 105.410 219.590 105.640 ;
        RECT 219.600 105.640 223.500 106.320 ;
        RECT 224.660 105.640 226.490 106.320 ;
        RECT 219.600 105.410 220.530 105.640 ;
        RECT 224.660 105.410 226.005 105.640 ;
        RECT 226.510 105.450 226.940 106.235 ;
        RECT 227.055 105.640 230.520 106.320 ;
        RECT 231.100 105.640 232.930 106.320 ;
        RECT 233.400 105.640 235.230 106.320 ;
        RECT 235.700 105.640 237.530 106.320 ;
        RECT 227.055 105.410 227.975 105.640 ;
        RECT 231.100 105.410 232.445 105.640 ;
        RECT 233.400 105.410 234.745 105.640 ;
        RECT 236.185 105.410 237.530 105.640 ;
        RECT 237.540 105.640 239.370 106.320 ;
        RECT 237.540 105.410 238.885 105.640 ;
        RECT 239.390 105.450 239.820 106.235 ;
        RECT 239.840 105.640 243.740 106.320 ;
        RECT 244.075 105.640 247.540 106.320 ;
        RECT 247.755 105.640 251.220 106.320 ;
        RECT 239.840 105.410 240.770 105.640 ;
        RECT 244.075 105.410 244.995 105.640 ;
        RECT 247.755 105.410 248.675 105.640 ;
        RECT 252.270 105.450 252.700 106.235 ;
        RECT 252.830 105.640 256.295 106.320 ;
        RECT 255.375 105.410 256.295 105.640 ;
        RECT 257.320 105.640 261.220 106.320 ;
        RECT 261.460 105.640 263.290 106.320 ;
        RECT 263.300 105.640 265.130 106.320 ;
        RECT 257.320 105.410 258.250 105.640 ;
        RECT 261.945 105.410 263.290 105.640 ;
        RECT 263.785 105.410 265.130 105.640 ;
        RECT 265.150 105.450 265.580 106.235 ;
        RECT 265.600 105.640 267.430 106.320 ;
        RECT 267.440 105.640 269.270 106.320 ;
        RECT 269.280 105.640 271.110 106.320 ;
        RECT 265.600 105.410 266.945 105.640 ;
        RECT 267.440 105.410 268.785 105.640 ;
        RECT 269.280 105.410 270.625 105.640 ;
        RECT 271.120 105.510 272.490 106.320 ;
        RECT 272.595 105.640 276.060 106.320 ;
        RECT 276.180 105.640 278.010 106.320 ;
        RECT 272.595 105.410 273.515 105.640 ;
        RECT 276.180 105.410 277.525 105.640 ;
        RECT 278.030 105.450 278.460 106.235 ;
        RECT 278.480 105.640 287.670 106.320 ;
        RECT 287.680 105.640 289.510 106.320 ;
        RECT 278.480 105.410 279.400 105.640 ;
        RECT 282.230 105.420 283.160 105.640 ;
        RECT 287.680 105.410 289.025 105.640 ;
        RECT 289.520 105.510 290.890 106.320 ;
        RECT 290.910 105.450 291.340 106.235 ;
        RECT 291.360 105.640 293.190 106.320 ;
        RECT 291.360 105.410 292.705 105.640 ;
        RECT 293.200 105.510 294.570 106.320 ;
        RECT 294.580 105.640 303.770 106.320 ;
        RECT 299.090 105.420 300.020 105.640 ;
        RECT 302.850 105.410 303.770 105.640 ;
        RECT 303.790 105.450 304.220 106.235 ;
        RECT 304.240 105.640 306.070 106.320 ;
        RECT 307.000 105.640 308.830 106.320 ;
        RECT 304.240 105.410 305.585 105.640 ;
        RECT 307.485 105.410 308.830 105.640 ;
        RECT 309.760 105.510 311.130 106.320 ;
      LAYER nwell ;
        RECT 161.905 102.290 311.325 105.120 ;
      LAYER pwell ;
        RECT 162.100 101.090 163.470 101.900 ;
        RECT 163.940 101.770 165.285 102.000 ;
        RECT 170.290 101.770 171.220 101.990 ;
        RECT 174.050 101.770 174.970 102.000 ;
        RECT 163.940 101.090 165.770 101.770 ;
        RECT 165.780 101.090 174.970 101.770 ;
        RECT 174.990 101.175 175.420 101.960 ;
        RECT 179.950 101.770 180.880 101.990 ;
        RECT 183.710 101.770 184.630 102.000 ;
        RECT 186.045 101.770 187.390 102.000 ;
        RECT 191.910 101.770 192.840 101.990 ;
        RECT 195.670 101.770 196.590 102.000 ;
        RECT 175.440 101.090 184.630 101.770 ;
        RECT 185.560 101.090 187.390 101.770 ;
        RECT 187.400 101.090 196.590 101.770 ;
        RECT 196.600 101.770 197.945 102.000 ;
        RECT 198.900 101.770 200.245 102.000 ;
        RECT 196.600 101.090 198.430 101.770 ;
        RECT 198.900 101.090 200.730 101.770 ;
        RECT 200.750 101.175 201.180 101.960 ;
        RECT 201.200 101.770 202.545 102.000 ;
        RECT 208.010 101.770 208.940 101.990 ;
        RECT 211.770 101.770 212.690 102.000 ;
        RECT 201.200 101.090 203.030 101.770 ;
        RECT 203.500 101.090 212.690 101.770 ;
        RECT 212.700 101.770 213.630 102.000 ;
        RECT 217.300 101.770 218.220 102.000 ;
        RECT 221.050 101.770 221.980 101.990 ;
        RECT 212.700 101.090 216.600 101.770 ;
        RECT 217.300 101.090 226.490 101.770 ;
        RECT 226.510 101.175 226.940 101.960 ;
        RECT 226.960 101.770 227.890 102.000 ;
        RECT 231.100 101.770 232.445 102.000 ;
        RECT 226.960 101.090 230.860 101.770 ;
        RECT 231.100 101.090 232.930 101.770 ;
        RECT 232.940 101.090 236.610 101.900 ;
        RECT 241.590 101.770 242.520 101.990 ;
        RECT 245.350 101.770 246.270 102.000 ;
        RECT 237.080 101.090 246.270 101.770 ;
        RECT 246.280 101.770 247.210 102.000 ;
        RECT 250.905 101.770 252.250 102.000 ;
        RECT 246.280 101.090 250.180 101.770 ;
        RECT 250.420 101.090 252.250 101.770 ;
        RECT 252.270 101.175 252.700 101.960 ;
        RECT 252.720 101.770 253.650 102.000 ;
        RECT 261.830 101.770 262.760 101.990 ;
        RECT 265.590 101.770 266.510 102.000 ;
        RECT 271.030 101.770 271.960 101.990 ;
        RECT 274.790 101.770 275.710 102.000 ;
        RECT 252.720 101.090 256.620 101.770 ;
        RECT 257.320 101.090 266.510 101.770 ;
        RECT 266.520 101.090 275.710 101.770 ;
        RECT 275.720 101.770 277.065 102.000 ;
        RECT 275.720 101.090 277.550 101.770 ;
        RECT 278.030 101.175 278.460 101.960 ;
        RECT 278.480 101.770 279.400 102.000 ;
        RECT 282.230 101.770 283.160 101.990 ;
        RECT 287.680 101.770 288.600 102.000 ;
        RECT 291.430 101.770 292.360 101.990 ;
        RECT 296.880 101.770 297.810 102.000 ;
        RECT 301.020 101.770 302.365 102.000 ;
        RECT 278.480 101.090 287.670 101.770 ;
        RECT 287.680 101.090 296.870 101.770 ;
        RECT 296.880 101.090 300.780 101.770 ;
        RECT 301.020 101.090 302.850 101.770 ;
        RECT 303.790 101.175 304.220 101.960 ;
        RECT 304.240 101.770 305.170 102.000 ;
        RECT 304.240 101.090 308.140 101.770 ;
        RECT 308.380 101.090 309.750 101.900 ;
        RECT 309.760 101.090 311.130 101.900 ;
        RECT 162.240 100.880 162.410 101.090 ;
        RECT 163.615 101.035 163.735 101.040 ;
        RECT 163.615 100.930 163.790 101.035 ;
        RECT 163.630 100.925 163.790 100.930 ;
        RECT 165.460 100.900 165.630 101.090 ;
        RECT 165.920 100.880 166.090 101.090 ;
        RECT 166.390 100.925 166.550 101.035 ;
        RECT 167.300 100.880 167.470 101.070 ;
        RECT 175.580 100.900 175.750 101.090 ;
        RECT 177.235 100.880 177.405 101.070 ;
        RECT 181.110 100.925 181.270 101.035 ;
        RECT 183.400 100.880 183.570 101.070 ;
        RECT 184.790 100.935 184.950 101.045 ;
        RECT 185.700 100.900 185.870 101.090 ;
        RECT 187.265 100.880 187.435 101.070 ;
        RECT 187.540 100.900 187.710 101.090 ;
        RECT 188.460 100.880 188.630 101.070 ;
        RECT 197.935 100.880 198.105 101.070 ;
        RECT 198.120 100.900 198.290 101.090 ;
        RECT 198.575 100.930 198.695 101.040 ;
        RECT 200.420 100.900 200.590 101.090 ;
        RECT 201.800 100.880 201.970 101.070 ;
        RECT 202.720 100.900 202.890 101.090 ;
        RECT 203.175 100.930 203.295 101.040 ;
        RECT 203.640 100.900 203.810 101.090 ;
        RECT 211.920 100.880 212.090 101.070 ;
        RECT 212.380 100.880 212.550 101.070 ;
        RECT 213.115 100.900 213.285 101.090 ;
        RECT 215.600 100.880 215.770 101.070 ;
        RECT 216.060 100.880 216.230 101.070 ;
        RECT 216.975 100.930 217.095 101.040 ;
        RECT 217.900 100.880 218.070 101.070 ;
        RECT 226.180 100.900 226.350 101.090 ;
        RECT 227.100 100.880 227.270 101.070 ;
        RECT 227.375 100.900 227.545 101.090 ;
        RECT 229.860 100.880 230.030 101.070 ;
        RECT 232.620 100.900 232.790 101.090 ;
        RECT 233.080 100.900 233.250 101.090 ;
        RECT 235.380 100.880 235.550 101.070 ;
        RECT 236.755 100.930 236.875 101.040 ;
        RECT 237.220 100.900 237.390 101.090 ;
        RECT 239.055 100.930 239.175 101.040 ;
        RECT 239.980 100.880 240.150 101.070 ;
        RECT 246.695 100.900 246.865 101.090 ;
        RECT 249.180 100.880 249.350 101.070 ;
        RECT 250.560 100.900 250.730 101.090 ;
        RECT 253.135 100.900 253.305 101.090 ;
        RECT 256.995 100.930 257.115 101.040 ;
        RECT 257.460 100.900 257.630 101.090 ;
        RECT 259.760 100.880 259.930 101.070 ;
        RECT 260.220 100.880 260.390 101.070 ;
        RECT 262.975 100.930 263.095 101.040 ;
        RECT 264.820 100.880 264.990 101.070 ;
        RECT 265.740 100.880 265.910 101.070 ;
        RECT 266.660 100.900 266.830 101.090 ;
        RECT 267.395 100.880 267.565 101.070 ;
        RECT 271.255 100.930 271.375 101.040 ;
        RECT 271.720 100.880 271.890 101.070 ;
        RECT 277.240 100.900 277.410 101.090 ;
        RECT 277.695 100.930 277.815 101.040 ;
        RECT 284.325 100.880 284.495 101.070 ;
        RECT 286.440 100.880 286.610 101.070 ;
        RECT 287.360 100.900 287.530 101.090 ;
        RECT 288.280 100.880 288.450 101.070 ;
        RECT 290.120 100.880 290.290 101.070 ;
        RECT 290.575 100.930 290.695 101.040 ;
        RECT 291.775 100.880 291.945 101.070 ;
        RECT 295.635 100.930 295.755 101.040 ;
        RECT 296.100 100.880 296.270 101.070 ;
        RECT 296.560 100.900 296.730 101.090 ;
        RECT 297.295 100.900 297.465 101.090 ;
        RECT 302.540 100.900 302.710 101.090 ;
        RECT 303.010 100.935 303.170 101.045 ;
        RECT 304.655 100.900 304.825 101.090 ;
        RECT 305.300 100.880 305.470 101.070 ;
        RECT 307.140 100.880 307.310 101.070 ;
        RECT 308.520 100.900 308.690 101.090 ;
        RECT 308.990 100.925 309.150 101.035 ;
        RECT 310.820 100.880 310.990 101.090 ;
        RECT 162.100 100.070 163.470 100.880 ;
        RECT 164.400 100.200 166.230 100.880 ;
        RECT 167.160 100.200 176.770 100.880 ;
        RECT 164.400 99.970 165.745 100.200 ;
        RECT 171.670 99.980 172.600 100.200 ;
        RECT 175.430 99.970 176.770 100.200 ;
        RECT 176.820 100.200 180.720 100.880 ;
        RECT 181.880 100.200 183.710 100.880 ;
        RECT 183.950 100.200 187.850 100.880 ;
        RECT 176.820 99.970 177.750 100.200 ;
        RECT 181.880 99.970 183.225 100.200 ;
        RECT 186.920 99.970 187.850 100.200 ;
        RECT 187.870 100.010 188.300 100.795 ;
        RECT 188.320 100.200 197.510 100.880 ;
        RECT 192.830 99.980 193.760 100.200 ;
        RECT 196.590 99.970 197.510 100.200 ;
        RECT 197.520 100.200 201.420 100.880 ;
        RECT 197.520 99.970 198.450 100.200 ;
        RECT 201.660 100.070 203.030 100.880 ;
        RECT 203.040 100.200 212.230 100.880 ;
        RECT 203.040 99.970 203.960 100.200 ;
        RECT 206.790 99.980 207.720 100.200 ;
        RECT 212.240 100.070 213.610 100.880 ;
        RECT 213.630 100.010 214.060 100.795 ;
        RECT 214.080 100.200 215.910 100.880 ;
        RECT 214.080 99.970 215.425 100.200 ;
        RECT 215.920 100.070 217.750 100.880 ;
        RECT 217.760 100.200 226.950 100.880 ;
        RECT 222.270 99.980 223.200 100.200 ;
        RECT 226.030 99.970 226.950 100.200 ;
        RECT 226.960 99.970 229.710 100.880 ;
        RECT 229.720 100.070 235.230 100.880 ;
        RECT 235.240 100.070 238.910 100.880 ;
        RECT 239.390 100.010 239.820 100.795 ;
        RECT 239.840 100.200 249.030 100.880 ;
        RECT 249.040 100.200 258.230 100.880 ;
        RECT 244.350 99.980 245.280 100.200 ;
        RECT 248.110 99.970 249.030 100.200 ;
        RECT 253.550 99.980 254.480 100.200 ;
        RECT 257.310 99.970 258.230 100.200 ;
        RECT 258.240 100.200 260.070 100.880 ;
        RECT 258.240 99.970 259.585 100.200 ;
        RECT 260.080 100.070 262.830 100.880 ;
        RECT 263.300 100.200 265.130 100.880 ;
        RECT 263.300 99.970 264.645 100.200 ;
        RECT 265.150 100.010 265.580 100.795 ;
        RECT 265.600 100.070 266.970 100.880 ;
        RECT 266.980 100.200 270.880 100.880 ;
        RECT 271.580 100.200 280.770 100.880 ;
        RECT 281.010 100.200 284.910 100.880 ;
        RECT 266.980 99.970 267.910 100.200 ;
        RECT 276.090 99.980 277.020 100.200 ;
        RECT 279.850 99.970 280.770 100.200 ;
        RECT 283.980 99.970 284.910 100.200 ;
        RECT 284.920 100.200 286.750 100.880 ;
        RECT 286.760 100.200 288.590 100.880 ;
        RECT 288.600 100.200 290.430 100.880 ;
        RECT 284.920 99.970 286.265 100.200 ;
        RECT 286.760 99.970 288.105 100.200 ;
        RECT 288.600 99.970 289.945 100.200 ;
        RECT 290.910 100.010 291.340 100.795 ;
        RECT 291.360 100.200 295.260 100.880 ;
        RECT 295.960 100.200 305.150 100.880 ;
        RECT 305.160 100.200 306.990 100.880 ;
        RECT 307.000 100.200 308.830 100.880 ;
        RECT 291.360 99.970 292.290 100.200 ;
        RECT 300.470 99.980 301.400 100.200 ;
        RECT 304.230 99.970 305.150 100.200 ;
        RECT 305.645 99.970 306.990 100.200 ;
        RECT 307.485 99.970 308.830 100.200 ;
        RECT 309.760 100.070 311.130 100.880 ;
      LAYER nwell ;
        RECT 161.905 96.850 311.325 99.680 ;
      LAYER pwell ;
        RECT 162.100 95.650 163.470 96.460 ;
        RECT 163.940 96.330 165.285 96.560 ;
        RECT 165.780 96.330 167.125 96.560 ;
        RECT 163.940 95.650 165.770 96.330 ;
        RECT 165.780 95.650 167.610 96.330 ;
        RECT 167.620 95.650 170.370 96.460 ;
        RECT 170.840 96.330 171.770 96.560 ;
        RECT 170.840 95.650 174.740 96.330 ;
        RECT 174.990 95.735 175.420 96.520 ;
        RECT 175.440 96.330 176.370 96.560 ;
        RECT 175.440 95.650 179.340 96.330 ;
        RECT 179.580 95.650 182.330 96.460 ;
        RECT 182.800 95.650 185.550 96.560 ;
        RECT 185.560 95.650 187.390 96.460 ;
        RECT 187.860 96.330 188.790 96.560 ;
        RECT 192.000 96.330 192.930 96.560 ;
        RECT 187.860 95.650 191.760 96.330 ;
        RECT 192.000 95.650 195.900 96.330 ;
        RECT 196.140 95.650 198.890 96.460 ;
        RECT 199.385 96.330 200.730 96.560 ;
        RECT 198.900 95.650 200.730 96.330 ;
        RECT 200.750 95.735 201.180 96.520 ;
        RECT 201.200 95.650 203.030 96.460 ;
        RECT 203.050 95.650 205.780 96.560 ;
        RECT 205.800 95.650 209.010 96.560 ;
        RECT 211.675 96.330 212.595 96.560 ;
        RECT 209.130 95.650 212.595 96.330 ;
        RECT 212.700 95.650 218.210 96.460 ;
        RECT 218.220 95.650 221.890 96.460 ;
        RECT 221.900 95.650 223.270 96.460 ;
        RECT 223.280 95.650 226.490 96.560 ;
        RECT 226.510 95.735 226.940 96.520 ;
        RECT 227.420 95.650 231.075 96.560 ;
        RECT 231.100 95.650 236.610 96.460 ;
        RECT 236.620 95.650 240.290 96.460 ;
        RECT 240.760 95.650 243.970 96.560 ;
        RECT 243.980 95.650 247.190 96.560 ;
        RECT 248.135 95.650 251.790 96.560 ;
        RECT 252.270 95.735 252.700 96.520 ;
        RECT 252.720 95.650 255.930 96.560 ;
        RECT 255.940 95.650 259.140 96.560 ;
        RECT 259.160 95.650 264.670 96.460 ;
        RECT 264.680 95.650 268.350 96.460 ;
        RECT 269.280 96.330 270.625 96.560 ;
        RECT 271.120 96.330 272.465 96.560 ;
        RECT 273.880 96.330 274.810 96.560 ;
        RECT 269.280 95.650 271.110 96.330 ;
        RECT 271.120 95.650 272.950 96.330 ;
        RECT 273.880 95.650 277.780 96.330 ;
        RECT 278.030 95.735 278.460 96.520 ;
        RECT 281.680 96.330 282.610 96.560 ;
        RECT 278.710 95.650 282.610 96.330 ;
        RECT 282.620 95.650 285.370 96.560 ;
        RECT 285.865 96.330 287.210 96.560 ;
        RECT 285.380 95.650 287.210 96.330 ;
        RECT 287.220 95.650 288.590 96.460 ;
        RECT 289.085 96.330 290.430 96.560 ;
        RECT 288.600 95.650 290.430 96.330 ;
        RECT 290.440 96.330 291.785 96.560 ;
        RECT 290.440 95.650 292.270 96.330 ;
        RECT 292.280 95.650 294.110 96.460 ;
        RECT 299.090 96.330 300.020 96.550 ;
        RECT 302.850 96.330 303.770 96.560 ;
        RECT 294.580 95.650 303.770 96.330 ;
        RECT 303.790 95.735 304.220 96.520 ;
        RECT 304.240 96.330 305.170 96.560 ;
        RECT 304.240 95.650 308.140 96.330 ;
        RECT 308.380 95.650 309.750 96.460 ;
        RECT 309.760 95.650 311.130 96.460 ;
        RECT 162.240 95.440 162.410 95.650 ;
        RECT 163.615 95.490 163.735 95.600 ;
        RECT 165.000 95.440 165.170 95.630 ;
        RECT 165.460 95.440 165.630 95.650 ;
        RECT 167.300 95.460 167.470 95.650 ;
        RECT 167.760 95.460 167.930 95.650 ;
        RECT 169.140 95.440 169.310 95.630 ;
        RECT 170.520 95.600 170.690 95.630 ;
        RECT 170.515 95.490 170.690 95.600 ;
        RECT 170.520 95.440 170.690 95.490 ;
        RECT 171.255 95.460 171.425 95.650 ;
        RECT 175.855 95.460 176.025 95.650 ;
        RECT 179.720 95.440 179.890 95.650 ;
        RECT 182.475 95.490 182.595 95.600 ;
        RECT 182.940 95.460 183.110 95.650 ;
        RECT 185.240 95.440 185.410 95.630 ;
        RECT 185.700 95.460 185.870 95.650 ;
        RECT 187.535 95.490 187.655 95.600 ;
        RECT 188.275 95.460 188.445 95.650 ;
        RECT 188.470 95.485 188.630 95.595 ;
        RECT 189.380 95.440 189.550 95.630 ;
        RECT 192.140 95.440 192.310 95.630 ;
        RECT 192.415 95.460 192.585 95.650 ;
        RECT 194.900 95.440 195.070 95.630 ;
        RECT 196.280 95.460 196.450 95.650 ;
        RECT 199.040 95.460 199.210 95.650 ;
        RECT 200.420 95.440 200.590 95.630 ;
        RECT 201.340 95.460 201.510 95.650 ;
        RECT 203.180 95.460 203.350 95.650 ;
        RECT 205.940 95.440 206.110 95.630 ;
        RECT 208.700 95.440 208.870 95.650 ;
        RECT 209.160 95.460 209.330 95.650 ;
        RECT 211.920 95.440 212.090 95.630 ;
        RECT 212.840 95.460 213.010 95.650 ;
        RECT 214.220 95.440 214.390 95.630 ;
        RECT 218.360 95.460 218.530 95.650 ;
        RECT 219.740 95.440 219.910 95.630 ;
        RECT 222.040 95.460 222.210 95.650 ;
        RECT 223.420 95.460 223.590 95.650 ;
        RECT 225.270 95.485 225.430 95.595 ;
        RECT 227.095 95.490 227.215 95.600 ;
        RECT 227.565 95.460 227.735 95.650 ;
        RECT 229.395 95.440 229.565 95.630 ;
        RECT 229.860 95.440 230.030 95.630 ;
        RECT 231.240 95.460 231.410 95.650 ;
        RECT 235.380 95.440 235.550 95.630 ;
        RECT 236.760 95.460 236.930 95.650 ;
        RECT 239.055 95.490 239.175 95.600 ;
        RECT 239.980 95.440 240.150 95.630 ;
        RECT 240.435 95.490 240.555 95.600 ;
        RECT 243.660 95.460 243.830 95.650 ;
        RECT 244.120 95.460 244.290 95.650 ;
        RECT 244.575 95.440 244.745 95.630 ;
        RECT 245.040 95.440 245.210 95.630 ;
        RECT 246.885 95.440 247.055 95.630 ;
        RECT 247.350 95.495 247.510 95.605 ;
        RECT 251.475 95.460 251.645 95.650 ;
        RECT 251.935 95.490 252.055 95.600 ;
        RECT 253.775 95.440 253.945 95.630 ;
        RECT 254.240 95.440 254.410 95.630 ;
        RECT 255.620 95.460 255.790 95.650 ;
        RECT 258.845 95.460 259.015 95.650 ;
        RECT 259.300 95.460 259.470 95.650 ;
        RECT 259.760 95.440 259.930 95.630 ;
        RECT 264.820 95.460 264.990 95.650 ;
        RECT 265.740 95.440 265.910 95.630 ;
        RECT 268.510 95.495 268.670 95.605 ;
        RECT 270.800 95.460 270.970 95.650 ;
        RECT 271.260 95.440 271.430 95.630 ;
        RECT 272.640 95.460 272.810 95.650 ;
        RECT 273.110 95.495 273.270 95.605 ;
        RECT 274.295 95.460 274.465 95.650 ;
        RECT 276.775 95.490 276.895 95.600 ;
        RECT 279.540 95.440 279.710 95.630 ;
        RECT 280.000 95.440 280.170 95.630 ;
        RECT 282.025 95.460 282.195 95.650 ;
        RECT 284.140 95.440 284.310 95.630 ;
        RECT 284.600 95.440 284.770 95.630 ;
        RECT 285.060 95.460 285.230 95.650 ;
        RECT 285.520 95.460 285.690 95.650 ;
        RECT 287.360 95.460 287.530 95.650 ;
        RECT 288.740 95.460 288.910 95.650 ;
        RECT 290.130 95.485 290.290 95.595 ;
        RECT 291.775 95.440 291.945 95.630 ;
        RECT 291.960 95.460 292.130 95.650 ;
        RECT 292.420 95.460 292.590 95.650 ;
        RECT 294.255 95.490 294.375 95.600 ;
        RECT 294.720 95.460 294.890 95.650 ;
        RECT 295.650 95.485 295.810 95.595 ;
        RECT 296.835 95.440 297.005 95.630 ;
        RECT 300.975 95.440 301.145 95.630 ;
        RECT 304.655 95.460 304.825 95.650 ;
        RECT 304.840 95.440 305.010 95.630 ;
        RECT 306.675 95.490 306.795 95.600 ;
        RECT 307.140 95.440 307.310 95.630 ;
        RECT 308.520 95.460 308.690 95.650 ;
        RECT 308.990 95.485 309.150 95.595 ;
        RECT 310.820 95.440 310.990 95.650 ;
        RECT 162.100 94.630 163.470 95.440 ;
        RECT 163.480 94.760 165.310 95.440 ;
        RECT 163.480 94.530 164.825 94.760 ;
        RECT 165.320 94.630 168.990 95.440 ;
        RECT 169.000 94.630 170.370 95.440 ;
        RECT 170.380 94.760 179.570 95.440 ;
        RECT 174.890 94.540 175.820 94.760 ;
        RECT 178.650 94.530 179.570 94.760 ;
        RECT 179.580 94.630 185.090 95.440 ;
        RECT 185.100 94.630 187.850 95.440 ;
        RECT 187.870 94.570 188.300 95.355 ;
        RECT 189.240 94.760 191.980 95.440 ;
        RECT 192.000 94.530 194.750 95.440 ;
        RECT 194.760 94.630 200.270 95.440 ;
        RECT 200.280 94.630 205.790 95.440 ;
        RECT 205.810 94.530 208.540 95.440 ;
        RECT 208.560 94.530 211.770 95.440 ;
        RECT 211.780 94.630 213.610 95.440 ;
        RECT 213.630 94.570 214.060 95.355 ;
        RECT 214.080 94.630 219.590 95.440 ;
        RECT 219.600 94.630 225.110 95.440 ;
        RECT 226.055 94.530 229.710 95.440 ;
        RECT 229.720 94.630 235.230 95.440 ;
        RECT 235.240 94.630 238.910 95.440 ;
        RECT 239.390 94.570 239.820 95.355 ;
        RECT 239.840 94.630 241.210 95.440 ;
        RECT 241.235 94.530 244.890 95.440 ;
        RECT 244.900 94.630 246.730 95.440 ;
        RECT 246.740 94.530 250.395 95.440 ;
        RECT 250.435 94.530 254.090 95.440 ;
        RECT 254.100 94.630 259.610 95.440 ;
        RECT 259.620 94.630 265.130 95.440 ;
        RECT 265.150 94.570 265.580 95.355 ;
        RECT 265.600 94.630 271.110 95.440 ;
        RECT 271.120 94.630 276.630 95.440 ;
        RECT 277.100 94.530 279.850 95.440 ;
        RECT 279.860 94.630 281.690 95.440 ;
        RECT 281.700 94.530 284.450 95.440 ;
        RECT 284.460 94.630 289.970 95.440 ;
        RECT 290.910 94.570 291.340 95.355 ;
        RECT 291.360 94.760 295.260 95.440 ;
        RECT 296.420 94.760 300.320 95.440 ;
        RECT 300.560 94.760 304.460 95.440 ;
        RECT 304.700 94.760 306.530 95.440 ;
        RECT 307.000 94.760 308.830 95.440 ;
        RECT 291.360 94.530 292.290 94.760 ;
        RECT 296.420 94.530 297.350 94.760 ;
        RECT 300.560 94.530 301.490 94.760 ;
        RECT 305.185 94.530 306.530 94.760 ;
        RECT 307.485 94.530 308.830 94.760 ;
        RECT 309.760 94.630 311.130 95.440 ;
      LAYER nwell ;
        RECT 161.905 91.410 311.325 94.240 ;
      LAYER pwell ;
        RECT 162.100 90.210 163.470 91.020 ;
        RECT 163.480 90.210 168.990 91.020 ;
        RECT 169.000 90.210 170.830 91.020 ;
        RECT 170.840 90.890 171.770 91.120 ;
        RECT 170.840 90.210 174.740 90.890 ;
        RECT 174.990 90.295 175.420 91.080 ;
        RECT 175.440 90.890 176.370 91.120 ;
        RECT 179.675 90.890 180.595 91.120 ;
        RECT 187.770 90.890 188.700 91.110 ;
        RECT 191.530 90.890 192.450 91.120 ;
        RECT 175.440 90.210 179.340 90.890 ;
        RECT 179.675 90.210 183.140 90.890 ;
        RECT 183.260 90.210 192.450 90.890 ;
        RECT 192.460 90.210 194.290 91.020 ;
        RECT 194.955 90.210 198.430 91.120 ;
        RECT 198.440 90.210 200.270 91.020 ;
        RECT 200.750 90.295 201.180 91.080 ;
        RECT 201.200 90.210 203.950 91.020 ;
        RECT 204.445 90.890 205.790 91.120 ;
        RECT 203.960 90.210 205.790 90.890 ;
        RECT 206.270 90.210 209.000 91.120 ;
        RECT 209.170 90.210 212.825 91.120 ;
        RECT 213.160 90.210 218.670 91.020 ;
        RECT 218.680 90.210 222.350 91.020 ;
        RECT 223.280 90.210 226.490 91.120 ;
        RECT 226.510 90.295 226.940 91.080 ;
        RECT 226.975 90.210 230.630 91.120 ;
        RECT 230.640 90.210 233.850 91.120 ;
        RECT 233.860 90.210 239.370 91.020 ;
        RECT 239.380 90.210 241.210 91.020 ;
        RECT 241.220 90.210 244.890 91.120 ;
        RECT 244.915 90.210 248.570 91.120 ;
        RECT 248.580 90.210 252.250 91.020 ;
        RECT 252.270 90.295 252.700 91.080 ;
        RECT 252.720 90.210 258.230 91.020 ;
        RECT 258.700 90.210 262.355 91.120 ;
        RECT 262.380 90.210 265.590 91.120 ;
        RECT 265.600 90.210 268.810 91.120 ;
        RECT 268.820 90.210 274.330 91.020 ;
        RECT 274.340 90.210 278.010 91.020 ;
        RECT 278.030 90.295 278.460 91.080 ;
        RECT 278.480 90.210 282.150 91.120 ;
        RECT 282.160 90.210 285.830 91.020 ;
        RECT 286.300 90.890 287.220 91.120 ;
        RECT 290.050 90.890 290.980 91.110 ;
        RECT 295.960 90.890 296.890 91.120 ;
        RECT 286.300 90.210 295.490 90.890 ;
        RECT 295.960 90.210 299.860 90.890 ;
        RECT 300.100 90.210 301.930 91.020 ;
        RECT 302.425 90.890 303.770 91.120 ;
        RECT 301.940 90.210 303.770 90.890 ;
        RECT 303.790 90.295 304.220 91.080 ;
        RECT 308.405 90.890 309.750 91.120 ;
        RECT 304.240 90.210 306.980 90.890 ;
        RECT 307.920 90.210 309.750 90.890 ;
        RECT 309.760 90.210 311.130 91.020 ;
        RECT 162.240 90.000 162.410 90.210 ;
        RECT 163.620 90.000 163.790 90.210 ;
        RECT 167.295 90.050 167.415 90.160 ;
        RECT 169.140 90.020 169.310 90.210 ;
        RECT 171.255 90.020 171.425 90.210 ;
        RECT 175.855 90.020 176.025 90.210 ;
        RECT 176.500 90.000 176.670 90.190 ;
        RECT 177.235 90.000 177.405 90.190 ;
        RECT 182.940 90.020 183.110 90.210 ;
        RECT 183.400 90.020 183.570 90.210 ;
        RECT 184.320 90.000 184.490 90.190 ;
        RECT 184.780 90.000 184.950 90.190 ;
        RECT 187.535 90.050 187.655 90.160 ;
        RECT 188.460 90.000 188.630 90.190 ;
        RECT 192.150 90.045 192.310 90.155 ;
        RECT 192.600 90.020 192.770 90.210 ;
        RECT 194.435 90.050 194.555 90.160 ;
        RECT 194.900 90.020 195.070 90.190 ;
        RECT 194.900 90.000 195.065 90.020 ;
        RECT 195.360 90.000 195.530 90.190 ;
        RECT 198.115 90.020 198.285 90.210 ;
        RECT 198.580 90.020 198.750 90.210 ;
        RECT 200.415 90.050 200.535 90.160 ;
        RECT 200.880 90.020 201.050 90.190 ;
        RECT 201.340 90.020 201.510 90.210 ;
        RECT 204.100 90.020 204.270 90.210 ;
        RECT 200.885 90.000 201.050 90.020 ;
        RECT 205.480 90.000 205.650 90.190 ;
        RECT 205.935 90.050 206.055 90.160 ;
        RECT 208.700 90.020 208.870 90.210 ;
        RECT 209.170 90.190 209.330 90.210 ;
        RECT 209.155 90.020 209.330 90.190 ;
        RECT 209.155 90.000 209.325 90.020 ;
        RECT 209.620 90.000 209.790 90.190 ;
        RECT 213.300 90.160 213.470 90.210 ;
        RECT 213.295 90.050 213.470 90.160 ;
        RECT 213.300 90.020 213.470 90.050 ;
        RECT 216.990 90.000 217.160 90.190 ;
        RECT 217.440 90.000 217.610 90.190 ;
        RECT 218.820 90.020 218.990 90.210 ;
        RECT 222.510 90.055 222.670 90.165 ;
        RECT 222.960 90.000 223.130 90.190 ;
        RECT 225.715 90.050 225.835 90.160 ;
        RECT 226.180 90.000 226.350 90.210 ;
        RECT 230.315 90.020 230.485 90.210 ;
        RECT 162.100 89.190 163.470 90.000 ;
        RECT 163.480 89.190 167.150 90.000 ;
        RECT 167.620 89.320 176.810 90.000 ;
        RECT 176.820 89.320 180.720 90.000 ;
        RECT 181.055 89.320 184.520 90.000 ;
        RECT 167.620 89.090 168.540 89.320 ;
        RECT 171.370 89.100 172.300 89.320 ;
        RECT 176.820 89.090 177.750 89.320 ;
        RECT 181.055 89.090 181.975 89.320 ;
        RECT 184.640 89.090 187.390 90.000 ;
        RECT 187.870 89.130 188.300 89.915 ;
        RECT 188.320 89.190 191.990 90.000 ;
        RECT 193.230 89.320 195.065 90.000 ;
        RECT 193.230 89.090 194.160 89.320 ;
        RECT 195.220 89.190 200.730 90.000 ;
        RECT 200.885 89.320 202.720 90.000 ;
        RECT 201.790 89.090 202.720 89.320 ;
        RECT 203.050 89.090 205.780 90.000 ;
        RECT 205.995 89.090 209.470 90.000 ;
        RECT 209.480 89.190 213.150 90.000 ;
        RECT 213.630 89.130 214.060 89.915 ;
        RECT 214.080 89.090 217.290 90.000 ;
        RECT 217.300 89.190 222.810 90.000 ;
        RECT 222.820 89.190 225.570 90.000 ;
        RECT 226.040 89.090 229.250 90.000 ;
        RECT 229.260 89.970 230.215 90.000 ;
        RECT 231.245 89.970 231.415 90.190 ;
        RECT 231.700 90.000 231.870 90.190 ;
        RECT 233.540 90.020 233.710 90.210 ;
        RECT 234.000 90.020 234.170 90.210 ;
        RECT 237.220 90.000 237.390 90.190 ;
        RECT 239.055 90.050 239.175 90.160 ;
        RECT 239.520 90.020 239.690 90.210 ;
        RECT 239.980 90.000 240.150 90.190 ;
        RECT 241.365 90.020 241.535 90.210 ;
        RECT 243.650 90.000 243.820 90.190 ;
        RECT 246.880 90.000 247.050 90.190 ;
        RECT 248.255 90.020 248.425 90.210 ;
        RECT 248.720 90.020 248.890 90.210 ;
        RECT 252.400 90.000 252.570 90.190 ;
        RECT 252.860 90.020 253.030 90.210 ;
        RECT 257.920 90.000 258.090 90.190 ;
        RECT 258.375 90.050 258.495 90.160 ;
        RECT 258.845 90.020 259.015 90.210 ;
        RECT 260.675 90.050 260.795 90.160 ;
        RECT 261.145 90.000 261.315 90.190 ;
        RECT 262.520 90.020 262.690 90.210 ;
        RECT 264.815 90.050 264.935 90.160 ;
        RECT 265.740 90.000 265.910 90.210 ;
        RECT 268.960 90.190 269.130 90.210 ;
        RECT 268.955 90.020 269.130 90.190 ;
        RECT 229.260 89.290 231.540 89.970 ;
        RECT 229.260 89.090 230.215 89.290 ;
        RECT 231.560 89.190 237.070 90.000 ;
        RECT 237.080 89.190 238.910 90.000 ;
        RECT 239.390 89.130 239.820 89.915 ;
        RECT 239.840 89.190 243.510 90.000 ;
        RECT 243.520 89.090 246.730 90.000 ;
        RECT 246.740 89.190 252.250 90.000 ;
        RECT 252.260 89.190 257.770 90.000 ;
        RECT 257.780 89.190 260.530 90.000 ;
        RECT 261.000 89.090 264.655 90.000 ;
        RECT 265.150 89.130 265.580 89.915 ;
        RECT 265.600 89.090 268.810 90.000 ;
        RECT 268.955 89.970 269.125 90.020 ;
        RECT 271.260 90.000 271.430 90.190 ;
        RECT 274.480 90.020 274.650 90.210 ;
        RECT 276.780 90.000 276.950 90.190 ;
        RECT 270.155 89.970 271.110 90.000 ;
        RECT 268.830 89.290 271.110 89.970 ;
        RECT 270.155 89.090 271.110 89.290 ;
        RECT 271.120 89.190 276.630 90.000 ;
        RECT 276.640 89.190 278.010 90.000 ;
        RECT 278.165 89.970 278.335 90.190 ;
        RECT 278.625 90.020 278.795 90.210 ;
        RECT 280.920 90.000 281.090 90.190 ;
        RECT 282.300 90.020 282.470 90.210 ;
        RECT 285.975 90.050 286.095 90.160 ;
        RECT 286.440 90.000 286.610 90.190 ;
        RECT 290.130 90.045 290.290 90.155 ;
        RECT 291.500 90.000 291.670 90.190 ;
        RECT 295.180 90.000 295.350 90.210 ;
        RECT 295.635 90.050 295.755 90.160 ;
        RECT 296.375 90.020 296.545 90.210 ;
        RECT 300.240 90.020 300.410 90.210 ;
        RECT 302.080 90.020 302.250 90.210 ;
        RECT 304.380 90.020 304.550 90.210 ;
        RECT 304.840 90.000 305.010 90.190 ;
        RECT 306.220 90.000 306.390 90.190 ;
        RECT 307.150 90.055 307.310 90.165 ;
        RECT 308.060 90.000 308.230 90.210 ;
        RECT 310.820 90.000 310.990 90.210 ;
        RECT 279.825 89.970 280.770 90.000 ;
        RECT 278.020 89.290 280.770 89.970 ;
        RECT 279.825 89.090 280.770 89.290 ;
        RECT 280.780 89.190 286.290 90.000 ;
        RECT 286.300 89.190 289.970 90.000 ;
        RECT 290.910 89.130 291.340 89.915 ;
        RECT 291.360 89.190 295.030 90.000 ;
        RECT 295.040 89.320 304.650 90.000 ;
        RECT 299.550 89.100 300.480 89.320 ;
        RECT 303.310 89.090 304.650 89.320 ;
        RECT 304.700 89.190 306.070 90.000 ;
        RECT 306.080 89.320 307.910 90.000 ;
        RECT 307.920 89.320 309.750 90.000 ;
        RECT 306.565 89.090 307.910 89.320 ;
        RECT 308.405 89.090 309.750 89.320 ;
        RECT 309.760 89.190 311.130 90.000 ;
      LAYER nwell ;
        RECT 161.905 85.970 311.325 88.800 ;
      LAYER pwell ;
        RECT 162.100 84.770 163.470 85.580 ;
        RECT 163.480 84.770 165.310 85.580 ;
        RECT 170.290 85.450 171.220 85.670 ;
        RECT 174.050 85.450 174.970 85.680 ;
        RECT 165.780 84.770 174.970 85.450 ;
        RECT 174.990 84.855 175.420 85.640 ;
        RECT 179.950 85.450 180.880 85.670 ;
        RECT 183.710 85.450 184.630 85.680 ;
        RECT 175.440 84.770 184.630 85.450 ;
        RECT 184.650 85.590 186.240 85.680 ;
        RECT 187.410 85.590 189.000 85.680 ;
        RECT 184.650 84.770 187.220 85.590 ;
        RECT 187.410 84.770 189.980 85.590 ;
        RECT 190.160 84.770 191.990 85.580 ;
        RECT 192.770 85.450 193.700 85.680 ;
        RECT 192.770 84.770 194.605 85.450 ;
        RECT 194.955 84.770 198.430 85.680 ;
        RECT 198.440 84.770 200.270 85.580 ;
        RECT 200.750 84.855 201.180 85.640 ;
        RECT 202.250 85.450 203.180 85.680 ;
        RECT 201.345 84.770 203.180 85.450 ;
        RECT 204.155 84.770 207.630 85.680 ;
        RECT 209.150 85.450 210.080 85.680 ;
        RECT 208.245 84.770 210.080 85.450 ;
        RECT 210.595 84.770 214.070 85.680 ;
        RECT 214.080 84.770 219.590 85.580 ;
        RECT 219.600 84.770 225.110 85.580 ;
        RECT 225.120 84.770 226.490 85.580 ;
        RECT 226.510 84.855 226.940 85.640 ;
        RECT 226.960 84.770 232.470 85.580 ;
        RECT 232.480 84.770 237.990 85.580 ;
        RECT 238.000 84.770 243.510 85.580 ;
        RECT 244.060 84.770 246.270 85.680 ;
        RECT 249.940 85.450 250.870 85.680 ;
        RECT 247.200 84.770 250.870 85.450 ;
        RECT 250.880 84.770 252.250 85.580 ;
        RECT 252.270 84.855 252.700 85.640 ;
        RECT 252.720 84.770 258.230 85.580 ;
        RECT 258.240 84.770 263.750 85.580 ;
        RECT 263.760 84.770 267.430 85.580 ;
        RECT 268.595 84.770 273.410 85.450 ;
        RECT 273.420 84.770 277.090 85.580 ;
        RECT 278.030 84.855 278.460 85.640 ;
        RECT 278.480 84.770 281.230 85.580 ;
        RECT 281.935 84.770 286.750 85.450 ;
        RECT 286.770 84.770 289.500 85.680 ;
        RECT 289.520 84.770 293.190 85.580 ;
        RECT 293.200 84.770 294.570 85.580 ;
        RECT 299.090 85.450 300.020 85.670 ;
        RECT 302.850 85.450 303.770 85.680 ;
        RECT 294.580 84.770 303.770 85.450 ;
        RECT 303.790 84.855 304.220 85.640 ;
        RECT 304.240 84.770 306.070 85.580 ;
        RECT 306.540 84.770 307.910 85.550 ;
        RECT 308.405 85.450 309.750 85.680 ;
        RECT 307.920 84.770 309.750 85.450 ;
        RECT 309.760 84.770 311.130 85.580 ;
        RECT 162.240 84.560 162.410 84.770 ;
        RECT 163.620 84.560 163.790 84.770 ;
        RECT 165.455 84.610 165.575 84.720 ;
        RECT 165.920 84.580 166.090 84.770 ;
        RECT 166.375 84.610 166.495 84.720 ;
        RECT 166.840 84.560 167.010 84.750 ;
        RECT 175.580 84.580 175.750 84.770 ;
        RECT 187.080 84.750 187.220 84.770 ;
        RECT 189.840 84.750 189.980 84.770 ;
        RECT 176.040 84.560 176.210 84.750 ;
        RECT 181.560 84.560 181.730 84.750 ;
        RECT 186.620 84.580 186.790 84.750 ;
        RECT 187.080 84.580 187.250 84.750 ;
        RECT 189.840 84.580 190.010 84.750 ;
        RECT 190.300 84.580 190.470 84.770 ;
        RECT 194.440 84.750 194.605 84.770 ;
        RECT 190.760 84.580 190.930 84.750 ;
        RECT 186.620 84.560 186.760 84.580 ;
        RECT 190.760 84.560 190.900 84.580 ;
        RECT 191.220 84.560 191.390 84.750 ;
        RECT 192.135 84.610 192.255 84.720 ;
        RECT 193.060 84.560 193.230 84.750 ;
        RECT 194.440 84.580 194.610 84.750 ;
        RECT 198.115 84.580 198.285 84.770 ;
        RECT 198.580 84.580 198.750 84.770 ;
        RECT 201.345 84.750 201.510 84.770 ;
        RECT 200.420 84.720 200.590 84.750 ;
        RECT 200.415 84.610 200.590 84.720 ;
        RECT 200.420 84.560 200.590 84.610 ;
        RECT 200.880 84.560 201.050 84.750 ;
        RECT 201.340 84.580 201.510 84.750 ;
        RECT 203.635 84.610 203.755 84.720 ;
        RECT 204.560 84.560 204.730 84.750 ;
        RECT 205.940 84.560 206.110 84.750 ;
        RECT 207.315 84.580 207.485 84.770 ;
        RECT 208.245 84.750 208.410 84.770 ;
        RECT 207.775 84.610 207.895 84.720 ;
        RECT 208.240 84.580 208.410 84.750 ;
        RECT 208.700 84.560 208.870 84.750 ;
        RECT 213.755 84.580 213.925 84.770 ;
        RECT 214.220 84.580 214.390 84.770 ;
        RECT 217.435 84.560 217.605 84.750 ;
        RECT 217.900 84.560 218.070 84.750 ;
        RECT 219.740 84.580 219.910 84.770 ;
        RECT 223.420 84.560 223.590 84.750 ;
        RECT 225.260 84.580 225.430 84.770 ;
        RECT 227.100 84.560 227.270 84.770 ;
        RECT 230.320 84.560 230.490 84.750 ;
        RECT 232.620 84.580 232.790 84.770 ;
        RECT 235.840 84.560 236.010 84.750 ;
        RECT 238.140 84.580 238.310 84.770 ;
        RECT 239.990 84.605 240.150 84.715 ;
        RECT 242.275 84.560 242.445 84.750 ;
        RECT 243.655 84.610 243.775 84.720 ;
        RECT 245.955 84.560 246.125 84.770 ;
        RECT 246.430 84.615 246.590 84.725 ;
        RECT 247.340 84.580 247.510 84.770 ;
        RECT 248.260 84.580 248.430 84.750 ;
        RECT 248.260 84.560 248.410 84.580 ;
        RECT 248.720 84.560 248.890 84.750 ;
        RECT 250.560 84.560 250.730 84.750 ;
        RECT 251.020 84.580 251.190 84.770 ;
        RECT 252.860 84.580 253.030 84.770 ;
        RECT 253.780 84.560 253.950 84.750 ;
        RECT 254.240 84.560 254.410 84.750 ;
        RECT 258.380 84.580 258.550 84.770 ;
        RECT 259.770 84.605 259.930 84.715 ;
        RECT 162.100 83.750 163.470 84.560 ;
        RECT 163.480 83.750 166.230 84.560 ;
        RECT 166.700 83.880 175.890 84.560 ;
        RECT 171.210 83.660 172.140 83.880 ;
        RECT 174.970 83.650 175.890 83.880 ;
        RECT 175.900 83.750 181.410 84.560 ;
        RECT 181.420 83.750 184.170 84.560 ;
        RECT 184.190 83.740 186.760 84.560 ;
        RECT 184.190 83.650 185.780 83.740 ;
        RECT 187.870 83.690 188.300 84.475 ;
        RECT 188.330 83.740 190.900 84.560 ;
        RECT 191.080 83.750 192.910 84.560 ;
        RECT 192.920 83.750 195.010 84.560 ;
        RECT 195.915 83.880 200.730 84.560 ;
        RECT 200.740 83.750 204.410 84.560 ;
        RECT 204.420 83.750 205.790 84.560 ;
        RECT 205.800 83.750 207.890 84.560 ;
        RECT 208.560 83.880 213.375 84.560 ;
        RECT 188.330 83.650 189.920 83.740 ;
        RECT 213.630 83.690 214.060 84.475 ;
        RECT 214.275 83.650 217.750 84.560 ;
        RECT 217.760 83.750 223.270 84.560 ;
        RECT 223.280 83.750 226.950 84.560 ;
        RECT 226.960 83.650 230.170 84.560 ;
        RECT 230.180 83.750 235.690 84.560 ;
        RECT 235.700 83.750 239.370 84.560 ;
        RECT 239.390 83.690 239.820 84.475 ;
        RECT 240.820 83.650 242.590 84.560 ;
        RECT 242.615 83.650 246.270 84.560 ;
        RECT 246.480 83.740 248.410 84.560 ;
        RECT 248.580 83.880 250.410 84.560 ;
        RECT 250.420 83.880 252.250 84.560 ;
        RECT 252.260 83.880 254.090 84.560 ;
        RECT 246.480 83.650 247.430 83.740 ;
        RECT 249.065 83.650 250.410 83.880 ;
        RECT 250.905 83.650 252.250 83.880 ;
        RECT 254.100 83.750 259.610 84.560 ;
        RECT 260.685 84.530 260.855 84.750 ;
        RECT 263.440 84.560 263.610 84.750 ;
        RECT 263.900 84.580 264.070 84.770 ;
        RECT 265.740 84.580 265.910 84.750 ;
        RECT 267.590 84.615 267.750 84.725 ;
        RECT 268.035 84.610 268.155 84.720 ;
        RECT 265.760 84.560 265.910 84.580 ;
        RECT 271.260 84.560 271.430 84.750 ;
        RECT 271.720 84.560 271.890 84.750 ;
        RECT 273.100 84.580 273.270 84.770 ;
        RECT 273.560 84.580 273.730 84.770 ;
        RECT 277.240 84.580 277.410 84.750 ;
        RECT 278.620 84.580 278.790 84.770 ;
        RECT 277.270 84.560 277.410 84.580 ;
        RECT 280.000 84.560 280.170 84.750 ;
        RECT 281.375 84.610 281.495 84.720 ;
        RECT 284.600 84.560 284.770 84.750 ;
        RECT 285.060 84.560 285.230 84.750 ;
        RECT 286.440 84.580 286.610 84.770 ;
        RECT 286.900 84.580 287.070 84.770 ;
        RECT 289.660 84.580 289.830 84.770 ;
        RECT 290.575 84.610 290.695 84.720 ;
        RECT 293.340 84.580 293.510 84.770 ;
        RECT 293.800 84.560 293.970 84.750 ;
        RECT 294.260 84.560 294.430 84.750 ;
        RECT 294.720 84.580 294.890 84.770 ;
        RECT 296.100 84.560 296.270 84.750 ;
        RECT 304.380 84.580 304.550 84.770 ;
        RECT 305.300 84.560 305.470 84.750 ;
        RECT 306.215 84.610 306.335 84.720 ;
        RECT 307.600 84.580 307.770 84.770 ;
        RECT 308.060 84.580 308.230 84.770 ;
        RECT 308.990 84.605 309.150 84.715 ;
        RECT 310.820 84.560 310.990 84.770 ;
        RECT 262.345 84.530 263.290 84.560 ;
        RECT 260.540 83.850 263.290 84.530 ;
        RECT 262.345 83.650 263.290 83.850 ;
        RECT 263.300 83.750 265.130 84.560 ;
        RECT 265.150 83.690 265.580 84.475 ;
        RECT 265.760 83.740 267.690 84.560 ;
        RECT 266.740 83.650 267.690 83.740 ;
        RECT 268.360 83.650 271.520 84.560 ;
        RECT 271.580 83.750 277.090 84.560 ;
        RECT 277.270 83.740 279.840 84.560 ;
        RECT 279.860 83.750 281.690 84.560 ;
        RECT 278.250 83.650 279.840 83.740 ;
        RECT 281.700 83.650 284.860 84.560 ;
        RECT 284.920 83.750 290.430 84.560 ;
        RECT 290.910 83.690 291.340 84.475 ;
        RECT 292.020 83.750 294.110 84.560 ;
        RECT 294.120 83.750 295.950 84.560 ;
        RECT 295.960 83.880 305.150 84.560 ;
        RECT 300.470 83.660 301.400 83.880 ;
        RECT 304.230 83.650 305.150 83.880 ;
        RECT 305.160 83.750 308.830 84.560 ;
        RECT 309.760 83.750 311.130 84.560 ;
      LAYER nwell ;
        RECT 161.905 80.530 311.325 83.360 ;
      LAYER pwell ;
        RECT 162.100 79.330 163.470 80.140 ;
        RECT 163.480 79.330 168.990 80.140 ;
        RECT 169.000 79.330 170.830 80.140 ;
        RECT 170.840 80.010 171.770 80.240 ;
        RECT 170.840 79.330 174.740 80.010 ;
        RECT 174.990 79.415 175.420 80.200 ;
        RECT 175.440 80.010 176.370 80.240 ;
        RECT 175.440 79.330 179.340 80.010 ;
        RECT 179.580 79.330 185.090 80.140 ;
        RECT 185.100 79.330 188.770 80.140 ;
        RECT 188.780 79.330 191.940 80.240 ;
        RECT 192.000 79.330 193.830 80.140 ;
        RECT 194.300 79.330 197.050 80.240 ;
        RECT 197.060 79.330 200.730 80.140 ;
        RECT 200.750 79.415 201.180 80.200 ;
        RECT 201.200 79.330 204.870 80.140 ;
        RECT 204.880 79.330 211.390 80.240 ;
        RECT 211.780 79.330 218.290 80.240 ;
        RECT 218.680 79.330 222.350 80.140 ;
        RECT 222.360 79.330 223.730 80.140 ;
        RECT 225.080 80.040 226.490 80.240 ;
        RECT 223.755 79.360 226.490 80.040 ;
        RECT 226.510 79.415 226.940 80.200 ;
        RECT 162.240 79.120 162.410 79.330 ;
        RECT 163.620 79.120 163.790 79.330 ;
        RECT 169.140 79.140 169.310 79.330 ;
        RECT 170.060 79.120 170.230 79.310 ;
        RECT 171.255 79.140 171.425 79.330 ;
        RECT 175.855 79.140 176.025 79.330 ;
        RECT 179.720 79.140 179.890 79.330 ;
        RECT 179.995 79.120 180.165 79.310 ;
        RECT 183.870 79.165 184.030 79.275 ;
        RECT 184.775 79.120 184.945 79.310 ;
        RECT 185.240 79.140 185.410 79.330 ;
        RECT 188.455 79.170 188.575 79.280 ;
        RECT 191.680 79.140 191.850 79.330 ;
        RECT 192.140 79.140 192.310 79.330 ;
        RECT 193.520 79.120 193.690 79.310 ;
        RECT 193.980 79.280 194.150 79.310 ;
        RECT 193.975 79.170 194.150 79.280 ;
        RECT 162.100 78.310 163.470 79.120 ;
        RECT 163.480 78.310 168.990 79.120 ;
        RECT 169.920 78.440 179.530 79.120 ;
        RECT 174.430 78.220 175.360 78.440 ;
        RECT 178.190 78.210 179.530 78.440 ;
        RECT 179.580 78.440 183.480 79.120 ;
        RECT 179.580 78.210 180.510 78.440 ;
        RECT 184.650 78.210 187.850 79.120 ;
        RECT 187.870 78.250 188.300 79.035 ;
        RECT 189.015 78.440 193.830 79.120 ;
        RECT 193.980 79.090 194.150 79.170 ;
        RECT 196.740 79.140 196.910 79.330 ;
        RECT 197.200 79.140 197.370 79.330 ;
        RECT 199.955 79.120 200.125 79.310 ;
        RECT 200.420 79.120 200.590 79.310 ;
        RECT 201.340 79.140 201.510 79.330 ;
        RECT 204.095 79.170 204.215 79.280 ;
        RECT 195.180 79.090 196.560 79.120 ;
        RECT 193.855 78.410 196.560 79.090 ;
        RECT 195.180 78.210 196.560 78.410 ;
        RECT 196.795 78.210 200.270 79.120 ;
        RECT 200.280 78.310 203.950 79.120 ;
        RECT 204.560 79.090 204.730 79.310 ;
        RECT 205.025 79.140 205.195 79.330 ;
        RECT 208.240 79.120 208.410 79.310 ;
        RECT 211.000 79.140 211.170 79.310 ;
        RECT 211.925 79.140 212.095 79.330 ;
        RECT 213.295 79.170 213.415 79.280 ;
        RECT 211.005 79.120 211.170 79.140 ;
        RECT 214.220 79.120 214.390 79.310 ;
        RECT 218.820 79.140 218.990 79.330 ;
        RECT 219.740 79.120 219.910 79.310 ;
        RECT 222.500 79.140 222.670 79.330 ;
        RECT 223.415 79.170 223.535 79.280 ;
        RECT 223.880 79.120 224.050 79.360 ;
        RECT 225.095 79.330 226.490 79.360 ;
        RECT 226.960 79.330 228.790 80.140 ;
        RECT 228.815 79.330 232.470 80.240 ;
        RECT 232.490 79.330 235.220 80.240 ;
        RECT 235.240 79.330 238.910 80.140 ;
        RECT 239.380 79.330 242.590 80.240 ;
        RECT 242.600 79.330 246.255 80.240 ;
        RECT 246.280 80.040 247.665 80.240 ;
        RECT 246.280 79.360 249.950 80.040 ;
        RECT 246.280 79.330 247.650 79.360 ;
        RECT 226.635 79.170 226.755 79.280 ;
        RECT 206.720 79.090 208.090 79.120 ;
        RECT 204.420 78.410 208.090 79.090 ;
        RECT 206.705 78.210 208.090 78.410 ;
        RECT 208.100 78.310 210.850 79.120 ;
        RECT 211.005 78.440 212.840 79.120 ;
        RECT 211.910 78.210 212.840 78.440 ;
        RECT 213.630 78.250 214.060 79.035 ;
        RECT 214.080 78.310 219.590 79.120 ;
        RECT 219.600 78.310 223.270 79.120 ;
        RECT 223.740 78.210 226.490 79.120 ;
        RECT 227.100 79.090 227.270 79.330 ;
        RECT 230.780 79.120 230.950 79.310 ;
        RECT 232.155 79.140 232.325 79.330 ;
        RECT 232.620 79.140 232.790 79.330 ;
        RECT 235.380 79.140 235.550 79.330 ;
        RECT 236.300 79.120 236.470 79.310 ;
        RECT 239.055 79.170 239.175 79.280 ;
        RECT 239.520 79.140 239.690 79.330 ;
        RECT 242.745 79.310 242.915 79.330 ;
        RECT 239.980 79.120 240.150 79.310 ;
        RECT 242.740 79.140 242.915 79.310 ;
        RECT 242.740 79.120 242.910 79.140 ;
        RECT 229.260 79.090 230.630 79.120 ;
        RECT 226.960 78.410 230.630 79.090 ;
        RECT 229.245 78.210 230.630 78.410 ;
        RECT 230.640 78.310 236.150 79.120 ;
        RECT 236.160 78.310 238.910 79.120 ;
        RECT 239.390 78.250 239.820 79.035 ;
        RECT 239.840 78.310 242.590 79.120 ;
        RECT 242.600 78.210 245.810 79.120 ;
        RECT 245.965 79.090 246.135 79.310 ;
        RECT 248.720 79.120 248.890 79.310 ;
        RECT 249.640 79.140 249.810 79.360 ;
        RECT 249.960 79.330 251.790 80.140 ;
        RECT 252.270 79.415 252.700 80.200 ;
        RECT 252.720 79.330 254.090 80.140 ;
        RECT 254.100 79.330 257.310 80.240 ;
        RECT 257.320 79.330 260.975 80.240 ;
        RECT 261.015 79.330 264.670 80.240 ;
        RECT 264.680 79.330 267.890 80.240 ;
        RECT 269.705 80.040 270.650 80.240 ;
        RECT 267.900 79.360 270.650 80.040 ;
        RECT 250.100 79.140 250.270 79.330 ;
        RECT 251.935 79.170 252.055 79.280 ;
        RECT 252.860 79.140 253.030 79.330 ;
        RECT 254.240 79.120 254.410 79.330 ;
        RECT 257.465 79.140 257.635 79.330 ;
        RECT 257.915 79.170 258.035 79.280 ;
        RECT 258.380 79.120 258.550 79.310 ;
        RECT 261.600 79.120 261.770 79.310 ;
        RECT 264.355 79.140 264.525 79.330 ;
        RECT 264.815 79.170 264.935 79.280 ;
        RECT 267.580 79.140 267.750 79.330 ;
        RECT 268.045 79.310 268.215 79.360 ;
        RECT 269.705 79.330 270.650 79.360 ;
        RECT 270.660 79.330 276.170 80.140 ;
        RECT 276.180 79.330 278.010 80.140 ;
        RECT 278.030 79.415 278.460 80.200 ;
        RECT 278.480 79.330 280.310 80.140 ;
        RECT 280.780 80.010 281.710 80.240 ;
        RECT 284.920 80.010 285.850 80.240 ;
        RECT 280.780 79.330 284.680 80.010 ;
        RECT 284.920 79.330 288.820 80.010 ;
        RECT 289.060 79.330 290.430 80.140 ;
        RECT 293.640 80.010 294.570 80.240 ;
        RECT 290.670 79.330 294.570 80.010 ;
        RECT 294.580 80.010 295.500 80.240 ;
        RECT 298.330 80.010 299.260 80.230 ;
        RECT 294.580 79.330 303.770 80.010 ;
        RECT 303.790 79.415 304.220 80.200 ;
        RECT 304.240 79.330 309.750 80.140 ;
        RECT 309.760 79.330 311.130 80.140 ;
        RECT 268.040 79.140 268.215 79.310 ;
        RECT 270.800 79.140 270.970 79.330 ;
        RECT 267.580 79.120 267.730 79.140 ;
        RECT 268.040 79.120 268.210 79.140 ;
        RECT 273.560 79.120 273.730 79.310 ;
        RECT 276.320 79.140 276.490 79.330 ;
        RECT 278.620 79.140 278.790 79.330 ;
        RECT 279.090 79.165 279.250 79.275 ;
        RECT 280.455 79.170 280.575 79.280 ;
        RECT 281.195 79.140 281.365 79.330 ;
        RECT 285.335 79.140 285.505 79.330 ;
        RECT 288.740 79.120 288.910 79.310 ;
        RECT 289.200 79.120 289.370 79.330 ;
        RECT 291.500 79.120 291.670 79.310 ;
        RECT 293.985 79.140 294.155 79.330 ;
        RECT 296.560 79.120 296.730 79.310 ;
        RECT 297.940 79.120 298.110 79.310 ;
        RECT 303.460 79.140 303.630 79.330 ;
        RECT 304.380 79.140 304.550 79.330 ;
        RECT 307.600 79.120 307.770 79.310 ;
        RECT 309.435 79.170 309.555 79.280 ;
        RECT 310.820 79.120 310.990 79.330 ;
        RECT 247.625 79.090 248.570 79.120 ;
        RECT 245.820 78.410 248.570 79.090 ;
        RECT 247.625 78.210 248.570 78.410 ;
        RECT 248.580 78.310 254.090 79.120 ;
        RECT 254.100 78.310 257.770 79.120 ;
        RECT 258.240 78.210 261.450 79.120 ;
        RECT 261.460 78.210 264.670 79.120 ;
        RECT 265.150 78.250 265.580 79.035 ;
        RECT 265.800 78.300 267.730 79.120 ;
        RECT 267.900 78.310 273.410 79.120 ;
        RECT 273.420 78.310 278.930 79.120 ;
        RECT 279.860 78.440 289.050 79.120 ;
        RECT 265.800 78.210 266.750 78.300 ;
        RECT 279.860 78.210 280.780 78.440 ;
        RECT 283.610 78.220 284.540 78.440 ;
        RECT 289.060 78.310 290.890 79.120 ;
        RECT 290.910 78.250 291.340 79.035 ;
        RECT 291.360 78.440 296.175 79.120 ;
        RECT 296.420 78.310 297.790 79.120 ;
        RECT 297.800 78.440 307.410 79.120 ;
        RECT 302.310 78.220 303.240 78.440 ;
        RECT 306.070 78.210 307.410 78.440 ;
        RECT 307.460 78.310 309.290 79.120 ;
        RECT 309.760 78.310 311.130 79.120 ;
      LAYER nwell ;
        RECT 161.905 75.090 311.325 77.920 ;
      LAYER pwell ;
        RECT 162.100 73.890 163.470 74.700 ;
        RECT 163.480 73.890 165.310 74.700 ;
        RECT 170.290 74.570 171.220 74.790 ;
        RECT 174.050 74.570 174.970 74.800 ;
        RECT 165.780 73.890 174.970 74.570 ;
        RECT 174.990 73.975 175.420 74.760 ;
        RECT 175.440 74.570 176.370 74.800 ;
        RECT 175.440 73.890 179.340 74.570 ;
        RECT 179.580 73.890 180.950 74.700 ;
        RECT 185.470 74.570 186.400 74.790 ;
        RECT 189.230 74.570 190.150 74.800 ;
        RECT 180.960 73.890 190.150 74.570 ;
        RECT 190.160 73.890 191.530 74.700 ;
        RECT 196.050 74.570 196.980 74.790 ;
        RECT 199.810 74.570 200.730 74.800 ;
        RECT 191.540 73.890 200.730 74.570 ;
        RECT 200.750 73.975 201.180 74.760 ;
        RECT 201.200 74.570 202.545 74.800 ;
        RECT 201.200 73.890 203.030 74.570 ;
        RECT 203.040 73.890 206.710 74.700 ;
        RECT 207.180 74.570 208.100 74.800 ;
        RECT 210.930 74.570 211.860 74.790 ;
        RECT 216.380 74.570 217.310 74.800 ;
        RECT 207.180 73.890 216.370 74.570 ;
        RECT 216.380 73.890 220.280 74.570 ;
        RECT 220.520 73.890 223.270 74.700 ;
        RECT 223.740 74.570 225.085 74.800 ;
        RECT 223.740 73.890 225.570 74.570 ;
        RECT 226.510 73.975 226.940 74.760 ;
        RECT 226.960 73.890 232.470 74.700 ;
        RECT 232.480 73.890 237.990 74.700 ;
        RECT 238.000 73.890 243.510 74.700 ;
        RECT 243.520 73.890 249.030 74.700 ;
        RECT 249.040 73.890 251.790 74.700 ;
        RECT 252.270 73.975 252.700 74.760 ;
        RECT 252.720 73.890 258.230 74.700 ;
        RECT 258.240 73.890 260.070 74.700 ;
        RECT 260.080 73.890 263.735 74.800 ;
        RECT 263.760 73.890 269.270 74.700 ;
        RECT 269.280 73.890 274.790 74.700 ;
        RECT 274.810 73.890 278.010 74.800 ;
        RECT 278.030 73.975 278.460 74.760 ;
        RECT 278.940 74.570 279.860 74.800 ;
        RECT 282.690 74.570 283.620 74.790 ;
        RECT 278.940 73.890 288.130 74.570 ;
        RECT 288.140 73.890 289.510 74.700 ;
        RECT 299.090 74.570 300.020 74.790 ;
        RECT 302.850 74.570 303.770 74.800 ;
        RECT 289.520 73.890 294.335 74.570 ;
        RECT 294.580 73.890 303.770 74.570 ;
        RECT 303.790 73.975 304.220 74.760 ;
        RECT 304.240 74.570 305.170 74.800 ;
        RECT 304.240 73.890 308.140 74.570 ;
        RECT 308.380 73.890 309.750 74.700 ;
        RECT 309.760 73.890 311.130 74.700 ;
        RECT 162.240 73.680 162.410 73.890 ;
        RECT 163.620 73.680 163.790 73.890 ;
        RECT 165.455 73.730 165.575 73.840 ;
        RECT 165.920 73.700 166.090 73.890 ;
        RECT 169.150 73.725 169.310 73.835 ;
        RECT 170.060 73.680 170.230 73.870 ;
        RECT 175.855 73.700 176.025 73.890 ;
        RECT 179.720 73.680 179.890 73.890 ;
        RECT 181.100 73.700 181.270 73.890 ;
        RECT 183.400 73.680 183.570 73.870 ;
        RECT 187.540 73.680 187.710 73.870 ;
        RECT 188.455 73.730 188.575 73.840 ;
        RECT 190.300 73.700 190.470 73.890 ;
        RECT 191.680 73.700 191.850 73.890 ;
        RECT 193.520 73.680 193.690 73.870 ;
        RECT 193.980 73.680 194.150 73.870 ;
        RECT 197.015 73.680 197.185 73.870 ;
        RECT 200.875 73.680 201.045 73.870 ;
        RECT 202.720 73.700 202.890 73.890 ;
        RECT 203.180 73.700 203.350 73.890 ;
        RECT 205.480 73.680 205.650 73.870 ;
        RECT 205.940 73.680 206.110 73.870 ;
        RECT 206.855 73.730 206.975 73.840 ;
        RECT 209.895 73.680 210.065 73.870 ;
        RECT 214.225 73.680 214.395 73.870 ;
        RECT 216.060 73.700 216.230 73.890 ;
        RECT 216.795 73.700 216.965 73.890 ;
        RECT 217.900 73.680 218.070 73.870 ;
        RECT 220.660 73.700 220.830 73.890 ;
        RECT 223.415 73.730 223.535 73.840 ;
        RECT 225.260 73.700 225.430 73.890 ;
        RECT 225.730 73.735 225.890 73.845 ;
        RECT 227.100 73.680 227.270 73.890 ;
        RECT 229.860 73.680 230.030 73.870 ;
        RECT 232.620 73.700 232.790 73.890 ;
        RECT 233.080 73.680 233.250 73.870 ;
        RECT 238.140 73.700 238.310 73.890 ;
        RECT 238.610 73.725 238.770 73.835 ;
        RECT 239.985 73.680 240.155 73.870 ;
        RECT 243.660 73.700 243.830 73.890 ;
        RECT 246.875 73.680 247.045 73.870 ;
        RECT 247.340 73.680 247.510 73.870 ;
        RECT 249.180 73.700 249.350 73.890 ;
        RECT 251.935 73.730 252.055 73.840 ;
        RECT 252.860 73.680 253.030 73.890 ;
        RECT 256.540 73.680 256.710 73.870 ;
        RECT 258.380 73.700 258.550 73.890 ;
        RECT 259.765 73.680 259.935 73.870 ;
        RECT 260.225 73.700 260.395 73.890 ;
        RECT 263.440 73.680 263.610 73.870 ;
        RECT 263.900 73.700 264.070 73.890 ;
        RECT 268.500 73.680 268.670 73.870 ;
        RECT 268.960 73.680 269.130 73.870 ;
        RECT 269.420 73.700 269.590 73.890 ;
        RECT 274.480 73.680 274.650 73.870 ;
        RECT 274.935 73.700 275.105 73.890 ;
        RECT 278.160 73.680 278.330 73.870 ;
        RECT 278.620 73.840 278.790 73.870 ;
        RECT 287.820 73.840 287.990 73.890 ;
        RECT 278.615 73.730 278.790 73.840 ;
        RECT 287.815 73.730 287.990 73.840 ;
        RECT 278.620 73.680 278.790 73.730 ;
        RECT 287.820 73.700 287.990 73.730 ;
        RECT 288.280 73.700 288.450 73.890 ;
        RECT 289.660 73.700 289.830 73.890 ;
        RECT 290.580 73.680 290.750 73.870 ;
        RECT 291.500 73.680 291.670 73.870 ;
        RECT 294.720 73.700 294.890 73.890 ;
        RECT 302.080 73.680 302.250 73.870 ;
        RECT 302.815 73.680 302.985 73.870 ;
        RECT 304.655 73.700 304.825 73.890 ;
        RECT 308.060 73.680 308.230 73.870 ;
        RECT 308.520 73.680 308.690 73.890 ;
        RECT 310.820 73.680 310.990 73.890 ;
        RECT 162.100 72.870 163.470 73.680 ;
        RECT 163.480 72.870 168.990 73.680 ;
        RECT 169.920 73.000 179.530 73.680 ;
        RECT 174.430 72.780 175.360 73.000 ;
        RECT 178.190 72.770 179.530 73.000 ;
        RECT 179.580 72.870 183.250 73.680 ;
        RECT 183.260 72.870 184.630 73.680 ;
        RECT 184.640 72.770 187.800 73.680 ;
        RECT 187.870 72.810 188.300 73.595 ;
        RECT 189.015 73.000 193.830 73.680 ;
        RECT 193.840 72.870 196.590 73.680 ;
        RECT 196.600 73.000 200.500 73.680 ;
        RECT 196.600 72.770 197.530 73.000 ;
        RECT 200.750 72.770 203.950 73.680 ;
        RECT 203.960 73.000 205.790 73.680 ;
        RECT 205.800 72.870 209.470 73.680 ;
        RECT 209.480 73.000 213.380 73.680 ;
        RECT 209.480 72.770 210.410 73.000 ;
        RECT 213.630 72.810 214.060 73.595 ;
        RECT 214.080 72.770 217.555 73.680 ;
        RECT 217.760 73.000 226.950 73.680 ;
        RECT 222.270 72.780 223.200 73.000 ;
        RECT 226.030 72.770 226.950 73.000 ;
        RECT 226.960 72.870 229.710 73.680 ;
        RECT 229.720 72.770 232.930 73.680 ;
        RECT 232.940 72.870 238.450 73.680 ;
        RECT 239.390 72.810 239.820 73.595 ;
        RECT 239.840 72.770 243.495 73.680 ;
        RECT 243.535 72.770 247.190 73.680 ;
        RECT 247.200 72.870 252.710 73.680 ;
        RECT 252.720 72.870 256.390 73.680 ;
        RECT 256.400 72.770 259.610 73.680 ;
        RECT 259.620 72.770 263.275 73.680 ;
        RECT 263.300 72.870 265.130 73.680 ;
        RECT 265.150 72.810 265.580 73.595 ;
        RECT 265.600 72.770 268.810 73.680 ;
        RECT 268.820 72.870 274.330 73.680 ;
        RECT 274.340 72.870 275.710 73.680 ;
        RECT 275.720 72.770 278.470 73.680 ;
        RECT 278.480 73.000 287.670 73.680 ;
        RECT 282.990 72.780 283.920 73.000 ;
        RECT 286.750 72.770 287.670 73.000 ;
        RECT 288.800 72.870 290.890 73.680 ;
        RECT 290.910 72.810 291.340 73.595 ;
        RECT 291.360 72.870 293.190 73.680 ;
        RECT 293.200 73.000 302.390 73.680 ;
        RECT 302.400 73.000 306.300 73.680 ;
        RECT 306.540 73.000 308.370 73.680 ;
        RECT 293.200 72.770 294.120 73.000 ;
        RECT 296.950 72.780 297.880 73.000 ;
        RECT 302.400 72.770 303.330 73.000 ;
        RECT 306.540 72.770 307.885 73.000 ;
        RECT 308.380 72.870 309.750 73.680 ;
        RECT 309.760 72.870 311.130 73.680 ;
      LAYER nwell ;
        RECT 161.905 69.650 311.325 72.480 ;
      LAYER pwell ;
        RECT 162.100 68.450 163.470 69.260 ;
        RECT 163.480 68.450 168.990 69.260 ;
        RECT 169.000 68.450 170.830 69.260 ;
        RECT 170.840 69.130 171.770 69.360 ;
        RECT 170.840 68.450 174.740 69.130 ;
        RECT 174.990 68.535 175.420 69.320 ;
        RECT 175.440 69.130 176.370 69.360 ;
        RECT 175.440 68.450 179.340 69.130 ;
        RECT 179.580 68.450 183.250 69.260 ;
        RECT 183.780 68.450 185.550 69.360 ;
        RECT 185.795 68.680 188.130 69.360 ;
        RECT 186.280 68.450 188.130 68.680 ;
        RECT 188.320 69.130 189.250 69.360 ;
        RECT 188.320 68.450 192.220 69.130 ;
        RECT 193.380 68.680 197.970 69.360 ;
        RECT 194.340 68.450 197.970 68.680 ;
        RECT 197.980 68.450 200.730 69.260 ;
        RECT 200.750 68.535 201.180 69.320 ;
        RECT 201.200 68.450 206.710 69.260 ;
        RECT 211.690 69.130 212.620 69.350 ;
        RECT 215.450 69.130 216.370 69.360 ;
        RECT 219.580 69.130 220.510 69.360 ;
        RECT 207.180 68.450 216.370 69.130 ;
        RECT 216.610 68.450 220.510 69.130 ;
        RECT 220.520 68.450 226.030 69.260 ;
        RECT 226.510 68.535 226.940 69.320 ;
        RECT 226.960 68.450 232.470 69.260 ;
        RECT 232.480 68.450 234.310 69.260 ;
        RECT 234.320 69.130 235.455 69.360 ;
        RECT 234.320 68.450 237.530 69.130 ;
        RECT 237.625 68.450 246.730 69.130 ;
        RECT 246.740 68.450 250.395 69.360 ;
        RECT 250.420 68.450 252.250 69.260 ;
        RECT 252.270 68.535 252.700 69.320 ;
        RECT 252.720 68.450 256.390 69.260 ;
        RECT 257.320 68.450 260.975 69.360 ;
        RECT 261.000 68.450 264.210 69.360 ;
        RECT 266.025 69.160 267.425 69.360 ;
        RECT 268.775 69.160 269.730 69.360 ;
        RECT 264.220 68.480 267.425 69.160 ;
        RECT 267.450 68.480 269.730 69.160 ;
        RECT 162.240 68.240 162.410 68.450 ;
        RECT 163.620 68.240 163.790 68.450 ;
        RECT 167.300 68.240 167.470 68.430 ;
        RECT 169.140 68.260 169.310 68.450 ;
        RECT 171.255 68.260 171.425 68.450 ;
        RECT 175.855 68.260 176.025 68.450 ;
        RECT 176.500 68.240 176.670 68.430 ;
        RECT 177.880 68.240 178.050 68.430 ;
        RECT 179.720 68.260 179.890 68.450 ;
        RECT 183.395 68.290 183.515 68.400 ;
        RECT 185.235 68.260 185.405 68.450 ;
        RECT 188.000 68.430 188.130 68.450 ;
        RECT 187.535 68.290 187.655 68.400 ;
        RECT 188.000 68.260 188.170 68.430 ;
        RECT 188.735 68.260 188.905 68.450 ;
        RECT 191.225 68.240 191.395 68.430 ;
        RECT 191.680 68.240 191.850 68.430 ;
        RECT 192.610 68.295 192.770 68.405 ;
        RECT 193.520 68.240 193.690 68.430 ;
        RECT 196.275 68.290 196.395 68.400 ;
        RECT 197.655 68.260 197.825 68.450 ;
        RECT 198.120 68.260 198.290 68.450 ;
        RECT 199.955 68.240 200.125 68.430 ;
        RECT 200.420 68.240 200.590 68.430 ;
        RECT 201.340 68.260 201.510 68.450 ;
        RECT 202.260 68.240 202.430 68.430 ;
        RECT 206.855 68.290 206.975 68.400 ;
        RECT 207.320 68.260 207.490 68.450 ;
        RECT 210.080 68.240 210.250 68.430 ;
        RECT 213.295 68.240 213.465 68.430 ;
        RECT 217.435 68.240 217.605 68.430 ;
        RECT 217.900 68.240 218.070 68.430 ;
        RECT 219.925 68.260 220.095 68.450 ;
        RECT 220.660 68.260 220.830 68.450 ;
        RECT 221.120 68.240 221.290 68.430 ;
        RECT 224.800 68.240 224.970 68.430 ;
        RECT 226.175 68.290 226.295 68.400 ;
        RECT 227.100 68.260 227.270 68.450 ;
        RECT 229.405 68.260 229.575 68.430 ;
        RECT 229.405 68.240 229.540 68.260 ;
        RECT 229.860 68.240 230.030 68.430 ;
        RECT 232.620 68.260 232.790 68.450 ;
        RECT 233.080 68.260 233.250 68.430 ;
        RECT 233.080 68.240 233.230 68.260 ;
        RECT 233.540 68.240 233.710 68.430 ;
        RECT 237.220 68.260 237.390 68.450 ;
        RECT 239.055 68.290 239.175 68.400 ;
        RECT 162.100 67.430 163.470 68.240 ;
        RECT 163.480 67.430 167.150 68.240 ;
        RECT 167.160 67.560 176.350 68.240 ;
        RECT 171.670 67.340 172.600 67.560 ;
        RECT 175.430 67.330 176.350 67.560 ;
        RECT 176.360 67.430 177.730 68.240 ;
        RECT 177.740 67.560 187.350 68.240 ;
        RECT 182.250 67.340 183.180 67.560 ;
        RECT 186.010 67.330 187.350 67.560 ;
        RECT 187.870 67.370 188.300 68.155 ;
        RECT 188.320 67.330 191.520 68.240 ;
        RECT 191.540 67.560 193.370 68.240 ;
        RECT 192.025 67.330 193.370 67.560 ;
        RECT 193.380 67.430 196.130 68.240 ;
        RECT 196.795 67.330 200.270 68.240 ;
        RECT 200.280 67.560 202.110 68.240 ;
        RECT 200.765 67.330 202.110 67.560 ;
        RECT 202.120 67.430 207.630 68.240 ;
        RECT 207.640 67.330 210.390 68.240 ;
        RECT 210.690 67.330 213.610 68.240 ;
        RECT 213.630 67.370 214.060 68.155 ;
        RECT 214.275 67.330 217.750 68.240 ;
        RECT 217.760 67.330 220.970 68.240 ;
        RECT 220.980 67.430 224.650 68.240 ;
        RECT 224.660 67.430 226.030 68.240 ;
        RECT 226.040 67.330 229.540 68.240 ;
        RECT 229.720 67.430 231.090 68.240 ;
        RECT 231.300 67.420 233.230 68.240 ;
        RECT 233.400 67.430 238.910 68.240 ;
        RECT 239.840 68.210 240.795 68.240 ;
        RECT 241.825 68.210 241.995 68.430 ;
        RECT 246.420 68.240 246.590 68.450 ;
        RECT 246.885 68.430 247.055 68.450 ;
        RECT 246.880 68.260 247.055 68.430 ;
        RECT 250.560 68.260 250.730 68.450 ;
        RECT 246.880 68.240 247.050 68.260 ;
        RECT 252.400 68.240 252.570 68.430 ;
        RECT 252.860 68.260 253.030 68.450 ;
        RECT 256.550 68.295 256.710 68.405 ;
        RECT 257.465 68.260 257.635 68.450 ;
        RECT 257.920 68.240 258.090 68.430 ;
        RECT 261.140 68.260 261.310 68.450 ;
        RECT 261.595 68.290 261.715 68.400 ;
        RECT 262.060 68.260 262.230 68.430 ;
        RECT 264.365 68.260 264.535 68.480 ;
        RECT 266.025 68.450 267.425 68.480 ;
        RECT 262.080 68.240 262.230 68.260 ;
        RECT 265.740 68.240 265.910 68.430 ;
        RECT 267.575 68.260 267.745 68.480 ;
        RECT 268.775 68.450 269.730 68.480 ;
        RECT 269.740 68.450 271.110 69.260 ;
        RECT 271.190 68.680 275.540 69.360 ;
        RECT 271.770 68.450 275.540 68.680 ;
        RECT 275.720 68.450 277.550 69.260 ;
        RECT 278.030 68.535 278.460 69.320 ;
        RECT 282.990 69.130 283.920 69.350 ;
        RECT 286.750 69.130 287.670 69.360 ;
        RECT 278.480 68.450 287.670 69.130 ;
        RECT 288.140 69.130 289.070 69.360 ;
        RECT 288.140 68.450 292.040 69.130 ;
        RECT 292.280 68.450 294.110 69.260 ;
        RECT 299.090 69.130 300.020 69.350 ;
        RECT 302.850 69.130 303.770 69.360 ;
        RECT 294.580 68.450 303.770 69.130 ;
        RECT 303.790 68.535 304.220 69.320 ;
        RECT 304.240 69.130 305.170 69.360 ;
        RECT 304.240 68.450 308.140 69.130 ;
        RECT 308.380 68.450 309.750 69.230 ;
        RECT 309.760 68.450 311.130 69.260 ;
        RECT 269.880 68.260 270.050 68.450 ;
        RECT 275.400 68.430 275.540 68.450 ;
        RECT 271.270 68.285 271.430 68.395 ;
        RECT 272.185 68.240 272.355 68.430 ;
        RECT 274.480 68.240 274.650 68.430 ;
        RECT 275.400 68.260 275.570 68.430 ;
        RECT 275.860 68.260 276.030 68.450 ;
        RECT 277.695 68.290 277.815 68.400 ;
        RECT 278.620 68.260 278.790 68.450 ;
        RECT 280.275 68.240 280.445 68.430 ;
        RECT 286.440 68.240 286.610 68.430 ;
        RECT 286.900 68.240 287.070 68.430 ;
        RECT 287.815 68.290 287.935 68.400 ;
        RECT 288.555 68.260 288.725 68.450 ;
        RECT 290.575 68.290 290.695 68.400 ;
        RECT 291.500 68.240 291.670 68.430 ;
        RECT 292.420 68.260 292.590 68.450 ;
        RECT 294.255 68.290 294.375 68.400 ;
        RECT 294.720 68.260 294.890 68.450 ;
        RECT 295.455 68.240 295.625 68.430 ;
        RECT 299.320 68.240 299.490 68.430 ;
        RECT 304.655 68.260 304.825 68.450 ;
        RECT 308.990 68.285 309.150 68.395 ;
        RECT 309.440 68.260 309.610 68.450 ;
        RECT 310.820 68.240 310.990 68.450 ;
        RECT 231.300 67.330 232.250 67.420 ;
        RECT 239.390 67.370 239.820 68.155 ;
        RECT 239.840 67.530 242.120 68.210 ;
        RECT 242.150 68.200 243.070 68.240 ;
        RECT 242.140 68.010 243.070 68.200 ;
        RECT 245.160 68.010 246.730 68.240 ;
        RECT 242.140 67.650 246.730 68.010 ;
        RECT 242.150 67.560 246.730 67.650 ;
        RECT 239.840 67.330 240.795 67.530 ;
        RECT 242.150 67.330 245.150 67.560 ;
        RECT 246.740 67.430 252.250 68.240 ;
        RECT 252.260 67.430 257.770 68.240 ;
        RECT 257.780 67.430 261.450 68.240 ;
        RECT 262.080 67.420 264.010 68.240 ;
        RECT 263.060 67.330 264.010 67.420 ;
        RECT 265.150 67.370 265.580 68.155 ;
        RECT 265.600 67.430 271.110 68.240 ;
        RECT 272.040 67.330 274.250 68.240 ;
        RECT 274.340 67.430 279.850 68.240 ;
        RECT 279.860 67.560 283.760 68.240 ;
        RECT 279.860 67.330 280.790 67.560 ;
        RECT 284.000 67.330 286.750 68.240 ;
        RECT 286.760 67.430 290.430 68.240 ;
        RECT 290.910 67.370 291.340 68.155 ;
        RECT 291.360 67.430 295.030 68.240 ;
        RECT 295.040 67.560 298.940 68.240 ;
        RECT 299.180 67.560 308.790 68.240 ;
        RECT 295.040 67.330 295.970 67.560 ;
        RECT 303.690 67.340 304.620 67.560 ;
        RECT 307.450 67.330 308.790 67.560 ;
        RECT 309.760 67.430 311.130 68.240 ;
      LAYER nwell ;
        RECT 161.905 64.210 311.325 67.040 ;
      LAYER pwell ;
        RECT 162.100 63.010 163.470 63.820 ;
        RECT 163.480 63.010 165.310 63.820 ;
        RECT 165.360 63.690 166.700 63.920 ;
        RECT 169.530 63.690 170.460 63.910 ;
        RECT 165.360 63.010 174.970 63.690 ;
        RECT 174.990 63.095 175.420 63.880 ;
        RECT 175.440 63.690 176.370 63.920 ;
        RECT 175.440 63.010 179.340 63.690 ;
        RECT 179.580 63.010 180.950 63.820 ;
        RECT 180.960 63.690 181.890 63.920 ;
        RECT 180.960 63.010 184.860 63.690 ;
        RECT 185.100 63.010 190.610 63.820 ;
        RECT 190.620 63.010 193.370 63.820 ;
        RECT 193.910 63.240 197.965 63.920 ;
        RECT 199.315 63.720 200.270 63.920 ;
        RECT 193.910 63.010 197.830 63.240 ;
        RECT 197.990 63.040 200.270 63.720 ;
        RECT 200.750 63.095 201.180 63.880 ;
        RECT 162.240 62.800 162.410 63.010 ;
        RECT 163.620 62.820 163.790 63.010 ;
        RECT 165.000 62.800 165.170 62.990 ;
        RECT 165.460 62.800 165.630 62.990 ;
        RECT 174.660 62.820 174.830 63.010 ;
        RECT 175.855 62.820 176.025 63.010 ;
        RECT 177.420 62.800 177.590 62.990 ;
        RECT 179.720 62.820 179.890 63.010 ;
        RECT 180.180 62.820 180.350 62.990 ;
        RECT 180.180 62.800 180.320 62.820 ;
        RECT 180.640 62.800 180.810 62.990 ;
        RECT 181.375 62.820 181.545 63.010 ;
        RECT 184.315 62.850 184.435 62.960 ;
        RECT 185.240 62.820 185.410 63.010 ;
        RECT 186.155 62.800 186.325 62.990 ;
        RECT 186.620 62.800 186.790 62.990 ;
        RECT 190.760 62.820 190.930 63.010 ;
        RECT 191.215 62.800 191.385 62.990 ;
        RECT 191.690 62.845 191.850 62.955 ;
        RECT 192.605 62.800 192.775 62.990 ;
        RECT 193.515 62.850 193.635 62.960 ;
        RECT 195.815 62.850 195.935 62.960 ;
        RECT 196.280 62.800 196.450 62.990 ;
        RECT 197.660 62.820 197.830 63.010 ;
        RECT 198.115 62.820 198.285 63.040 ;
        RECT 199.315 63.010 200.270 63.040 ;
        RECT 201.200 63.010 204.675 63.920 ;
        RECT 204.880 63.010 206.710 63.820 ;
        RECT 207.375 63.010 210.850 63.920 ;
        RECT 211.055 63.010 214.530 63.920 ;
        RECT 214.735 63.010 218.210 63.920 ;
        RECT 218.390 63.010 221.890 63.920 ;
        RECT 221.900 63.010 225.570 63.820 ;
        RECT 226.510 63.095 226.940 63.880 ;
        RECT 226.960 63.010 232.470 63.820 ;
        RECT 232.480 63.010 237.990 63.820 ;
        RECT 238.000 63.010 240.750 63.820 ;
        RECT 241.220 63.010 245.340 63.920 ;
        RECT 245.360 63.010 250.870 63.820 ;
        RECT 250.880 63.010 252.250 63.820 ;
        RECT 252.270 63.095 252.700 63.880 ;
        RECT 252.720 63.010 256.390 63.820 ;
        RECT 256.860 63.010 259.610 63.920 ;
        RECT 259.620 63.010 265.130 63.820 ;
        RECT 265.140 63.010 270.650 63.820 ;
        RECT 270.660 63.010 272.030 63.820 ;
        RECT 273.380 63.720 274.790 63.920 ;
        RECT 272.055 63.040 274.790 63.720 ;
        RECT 200.420 62.960 200.590 62.990 ;
        RECT 200.415 62.850 200.590 62.960 ;
        RECT 200.420 62.820 200.590 62.850 ;
        RECT 201.345 62.820 201.515 63.010 ;
        RECT 200.440 62.800 200.590 62.820 ;
        RECT 202.720 62.800 202.890 62.990 ;
        RECT 205.020 62.820 205.190 63.010 ;
        RECT 206.410 62.845 206.570 62.955 ;
        RECT 206.855 62.850 206.975 62.960 ;
        RECT 207.320 62.800 207.490 62.990 ;
        RECT 210.535 62.820 210.705 63.010 ;
        RECT 214.215 62.990 214.385 63.010 ;
        RECT 213.300 62.820 213.470 62.990 ;
        RECT 214.215 62.820 214.390 62.990 ;
        RECT 217.895 62.820 218.065 63.010 ;
        RECT 218.390 62.990 218.525 63.010 ;
        RECT 218.355 62.820 218.530 62.990 ;
        RECT 221.115 62.850 221.235 62.960 ;
        RECT 213.300 62.800 213.450 62.820 ;
        RECT 214.220 62.800 214.390 62.820 ;
        RECT 218.360 62.800 218.530 62.820 ;
        RECT 221.580 62.800 221.750 62.990 ;
        RECT 222.040 62.820 222.210 63.010 ;
        RECT 225.260 62.800 225.430 62.990 ;
        RECT 225.730 62.855 225.890 62.965 ;
        RECT 227.100 62.820 227.270 63.010 ;
        RECT 228.475 62.850 228.595 62.960 ;
        RECT 229.215 62.800 229.385 62.990 ;
        RECT 232.620 62.820 232.790 63.010 ;
        RECT 233.355 62.800 233.525 62.990 ;
        RECT 237.220 62.800 237.390 62.990 ;
        RECT 238.140 62.820 238.310 63.010 ;
        RECT 239.055 62.850 239.175 62.960 ;
        RECT 239.980 62.800 240.150 62.990 ;
        RECT 240.895 62.850 241.015 62.960 ;
        RECT 241.360 62.820 241.530 63.010 ;
        RECT 243.200 62.820 243.370 63.010 ;
        RECT 245.500 62.990 245.670 63.010 ;
        RECT 243.660 62.800 243.830 62.990 ;
        RECT 245.500 62.820 245.680 62.990 ;
        RECT 245.510 62.800 245.680 62.820 ;
        RECT 246.890 62.800 247.060 62.990 ;
        RECT 248.260 62.800 248.430 62.990 ;
        RECT 251.020 62.820 251.190 63.010 ;
        RECT 252.860 62.820 253.030 63.010 ;
        RECT 254.425 62.800 254.595 62.990 ;
        RECT 255.435 62.800 255.605 62.990 ;
        RECT 256.535 62.850 256.655 62.960 ;
        RECT 257.000 62.820 257.170 63.010 ;
        RECT 259.760 62.820 259.930 63.010 ;
        RECT 162.100 61.990 163.470 62.800 ;
        RECT 163.480 62.120 165.310 62.800 ;
        RECT 163.480 61.890 164.825 62.120 ;
        RECT 165.320 61.990 168.070 62.800 ;
        RECT 168.120 62.120 177.730 62.800 ;
        RECT 168.120 61.890 169.460 62.120 ;
        RECT 172.290 61.900 173.220 62.120 ;
        RECT 177.750 61.980 180.320 62.800 ;
        RECT 180.500 61.990 184.170 62.800 ;
        RECT 177.750 61.890 179.340 61.980 ;
        RECT 184.700 61.890 186.470 62.800 ;
        RECT 186.480 61.990 187.850 62.800 ;
        RECT 187.870 61.930 188.300 62.715 ;
        RECT 188.320 61.890 191.530 62.800 ;
        RECT 192.460 62.120 195.670 62.800 ;
        RECT 194.305 61.890 195.670 62.120 ;
        RECT 196.140 61.890 200.200 62.800 ;
        RECT 200.440 61.980 202.370 62.800 ;
        RECT 202.580 61.990 206.250 62.800 ;
        RECT 201.420 61.890 202.370 61.980 ;
        RECT 207.180 61.890 211.240 62.800 ;
        RECT 211.520 61.980 213.450 62.800 ;
        RECT 211.520 61.890 212.470 61.980 ;
        RECT 213.630 61.930 214.060 62.715 ;
        RECT 214.080 61.890 218.140 62.800 ;
        RECT 218.220 61.990 220.970 62.800 ;
        RECT 221.550 62.120 225.015 62.800 ;
        RECT 224.095 61.890 225.015 62.120 ;
        RECT 225.200 61.890 228.200 62.800 ;
        RECT 228.800 62.120 232.700 62.800 ;
        RECT 232.940 62.120 236.840 62.800 ;
        RECT 228.800 61.890 229.730 62.120 ;
        RECT 232.940 61.890 233.870 62.120 ;
        RECT 237.080 61.990 238.910 62.800 ;
        RECT 239.390 61.930 239.820 62.715 ;
        RECT 239.840 62.120 243.510 62.800 ;
        RECT 243.520 62.120 245.350 62.800 ;
        RECT 242.580 61.890 243.510 62.120 ;
        RECT 245.360 62.020 246.730 62.800 ;
        RECT 246.740 62.020 248.110 62.800 ;
        RECT 248.120 61.990 250.870 62.800 ;
        RECT 251.110 62.120 255.010 62.800 ;
        RECT 254.080 61.890 255.010 62.120 ;
        RECT 255.020 62.120 258.920 62.800 ;
        RECT 259.160 62.770 260.530 62.800 ;
        RECT 262.520 62.770 262.690 62.990 ;
        RECT 262.980 62.800 263.150 62.990 ;
        RECT 264.815 62.850 264.935 62.960 ;
        RECT 265.280 62.820 265.450 63.010 ;
        RECT 265.740 62.800 265.910 62.990 ;
        RECT 270.800 62.820 270.970 63.010 ;
        RECT 271.260 62.800 271.430 62.990 ;
        RECT 272.180 62.820 272.350 63.040 ;
        RECT 273.395 63.010 274.790 63.040 ;
        RECT 274.800 63.010 277.550 63.820 ;
        RECT 278.030 63.095 278.460 63.880 ;
        RECT 278.480 63.010 280.310 63.820 ;
        RECT 284.830 63.690 285.760 63.910 ;
        RECT 288.590 63.690 289.510 63.920 ;
        RECT 280.320 63.010 289.510 63.690 ;
        RECT 289.520 63.010 293.190 63.820 ;
        RECT 298.630 63.690 299.560 63.910 ;
        RECT 302.390 63.690 303.730 63.920 ;
        RECT 294.120 63.010 303.730 63.690 ;
        RECT 303.790 63.095 304.220 63.880 ;
        RECT 304.240 63.690 305.170 63.920 ;
        RECT 304.240 63.010 308.140 63.690 ;
        RECT 308.380 63.010 309.750 63.820 ;
        RECT 309.760 63.010 311.130 63.820 ;
        RECT 274.940 62.820 275.110 63.010 ;
        RECT 276.780 62.800 276.950 62.990 ;
        RECT 277.695 62.850 277.815 62.960 ;
        RECT 278.620 62.820 278.790 63.010 ;
        RECT 280.460 62.820 280.630 63.010 ;
        RECT 281.840 62.800 282.010 62.990 ;
        RECT 282.575 62.800 282.745 62.990 ;
        RECT 286.715 62.800 286.885 62.990 ;
        RECT 289.660 62.820 289.830 63.010 ;
        RECT 290.575 62.850 290.695 62.960 ;
        RECT 291.500 62.800 291.670 62.990 ;
        RECT 293.350 62.855 293.510 62.965 ;
        RECT 294.260 62.820 294.430 63.010 ;
        RECT 295.455 62.800 295.625 62.990 ;
        RECT 299.595 62.800 299.765 62.990 ;
        RECT 304.655 62.820 304.825 63.010 ;
        RECT 305.760 62.800 305.930 62.990 ;
        RECT 306.220 62.800 306.390 62.990 ;
        RECT 308.520 62.820 308.690 63.010 ;
        RECT 310.820 62.800 310.990 63.010 ;
        RECT 255.020 61.890 255.950 62.120 ;
        RECT 259.160 62.090 262.830 62.770 ;
        RECT 259.160 61.890 260.545 62.090 ;
        RECT 262.840 61.990 264.670 62.800 ;
        RECT 265.150 61.930 265.580 62.715 ;
        RECT 265.600 61.990 271.110 62.800 ;
        RECT 271.120 61.990 276.630 62.800 ;
        RECT 276.640 61.990 279.390 62.800 ;
        RECT 279.400 61.890 282.150 62.800 ;
        RECT 282.160 62.120 286.060 62.800 ;
        RECT 286.300 62.120 290.200 62.800 ;
        RECT 282.160 61.890 283.090 62.120 ;
        RECT 286.300 61.890 287.230 62.120 ;
        RECT 290.910 61.930 291.340 62.715 ;
        RECT 291.360 61.990 295.030 62.800 ;
        RECT 295.040 62.120 298.940 62.800 ;
        RECT 299.180 62.120 303.080 62.800 ;
        RECT 303.330 62.120 306.070 62.800 ;
        RECT 295.040 61.890 295.970 62.120 ;
        RECT 299.180 61.890 300.110 62.120 ;
        RECT 306.080 61.990 309.750 62.800 ;
        RECT 309.760 61.990 311.130 62.800 ;
      LAYER nwell ;
        RECT 161.905 58.770 311.325 61.600 ;
      LAYER pwell ;
        RECT 162.100 57.570 163.470 58.380 ;
        RECT 163.480 57.570 168.990 58.380 ;
        RECT 169.000 57.570 174.510 58.380 ;
        RECT 174.990 57.655 175.420 58.440 ;
        RECT 176.370 58.390 177.960 58.480 ;
        RECT 176.370 57.570 178.940 58.390 ;
        RECT 179.120 57.570 180.950 58.380 ;
        RECT 181.905 58.250 185.415 58.480 ;
        RECT 181.420 57.570 185.415 58.250 ;
        RECT 185.580 57.570 191.070 58.480 ;
        RECT 191.080 57.570 195.115 58.480 ;
        RECT 196.370 58.390 197.960 58.480 ;
        RECT 195.390 57.570 197.960 58.390 ;
        RECT 197.980 57.570 200.730 58.380 ;
        RECT 200.750 57.655 201.180 58.440 ;
        RECT 201.280 57.570 204.280 58.480 ;
        RECT 204.420 57.570 209.930 58.380 ;
        RECT 209.940 57.570 212.690 58.380 ;
        RECT 217.210 58.250 218.140 58.470 ;
        RECT 220.970 58.250 221.890 58.480 ;
        RECT 212.700 57.570 221.890 58.250 ;
        RECT 221.900 58.250 222.830 58.480 ;
        RECT 221.900 57.570 225.800 58.250 ;
        RECT 226.510 57.655 226.940 58.440 ;
        RECT 230.075 58.250 230.995 58.480 ;
        RECT 235.610 58.250 236.540 58.470 ;
        RECT 239.370 58.250 240.290 58.480 ;
        RECT 227.530 57.570 230.995 58.250 ;
        RECT 231.100 57.570 240.290 58.250 ;
        RECT 240.300 57.570 242.130 58.380 ;
        RECT 244.880 58.250 245.810 58.480 ;
        RECT 242.140 57.570 245.810 58.250 ;
        RECT 245.820 57.570 251.330 58.380 ;
        RECT 252.270 57.655 252.700 58.440 ;
        RECT 257.230 58.250 258.160 58.470 ;
        RECT 260.990 58.250 261.910 58.480 ;
        RECT 252.720 57.570 261.910 58.250 ;
        RECT 261.920 58.250 263.055 58.480 ;
        RECT 261.920 57.570 265.130 58.250 ;
        RECT 265.140 57.570 268.810 58.380 ;
        RECT 268.820 57.570 270.190 58.380 ;
        RECT 270.270 57.800 274.620 58.480 ;
        RECT 270.850 57.570 274.620 57.800 ;
        RECT 274.800 57.570 277.550 58.380 ;
        RECT 278.030 57.655 278.460 58.440 ;
        RECT 278.480 58.250 279.410 58.480 ;
        RECT 287.590 58.250 288.520 58.470 ;
        RECT 291.350 58.250 292.690 58.480 ;
        RECT 278.480 57.570 282.380 58.250 ;
        RECT 283.080 57.570 292.690 58.250 ;
        RECT 292.740 57.570 294.570 58.380 ;
        RECT 294.580 58.250 295.500 58.480 ;
        RECT 298.330 58.250 299.260 58.470 ;
        RECT 294.580 57.570 303.770 58.250 ;
        RECT 303.790 57.655 304.220 58.440 ;
        RECT 304.240 57.570 309.750 58.380 ;
        RECT 309.760 57.570 311.130 58.380 ;
        RECT 162.240 57.360 162.410 57.570 ;
        RECT 163.620 57.360 163.790 57.570 ;
        RECT 169.140 57.360 169.310 57.570 ;
        RECT 178.800 57.550 178.940 57.570 ;
        RECT 170.795 57.360 170.965 57.550 ;
        RECT 174.655 57.410 174.775 57.520 ;
        RECT 175.590 57.415 175.750 57.525 ;
        RECT 176.040 57.360 176.210 57.550 ;
        RECT 178.800 57.380 178.970 57.550 ;
        RECT 178.800 57.360 178.940 57.380 ;
        RECT 179.260 57.360 179.430 57.570 ;
        RECT 181.095 57.410 181.215 57.520 ;
        RECT 181.565 57.380 181.735 57.570 ;
        RECT 182.020 57.360 182.190 57.550 ;
        RECT 183.855 57.410 183.975 57.520 ;
        RECT 186.155 57.360 186.325 57.550 ;
        RECT 186.620 57.360 186.790 57.550 ;
        RECT 190.755 57.380 190.925 57.570 ;
        RECT 191.225 57.380 191.395 57.570 ;
        RECT 195.390 57.550 195.530 57.570 ;
        RECT 191.680 57.360 191.850 57.550 ;
        RECT 193.050 57.360 193.220 57.550 ;
        RECT 193.530 57.405 193.690 57.515 ;
        RECT 194.440 57.360 194.610 57.550 ;
        RECT 195.360 57.380 195.530 57.550 ;
        RECT 198.120 57.380 198.290 57.570 ;
        RECT 201.340 57.380 201.510 57.570 ;
        RECT 204.560 57.380 204.730 57.570 ;
        RECT 205.480 57.380 205.650 57.550 ;
        RECT 205.480 57.360 205.645 57.380 ;
        RECT 205.940 57.360 206.110 57.550 ;
        RECT 208.695 57.410 208.815 57.520 ;
        RECT 210.080 57.380 210.250 57.570 ;
        RECT 211.000 57.380 211.170 57.550 ;
        RECT 211.460 57.380 211.630 57.550 ;
        RECT 212.840 57.380 213.010 57.570 ;
        RECT 211.000 57.360 211.165 57.380 ;
        RECT 162.100 56.550 163.470 57.360 ;
        RECT 163.480 56.550 168.990 57.360 ;
        RECT 169.000 56.550 170.370 57.360 ;
        RECT 170.380 56.680 174.280 57.360 ;
        RECT 174.520 56.680 176.350 57.360 ;
        RECT 170.380 56.450 171.310 56.680 ;
        RECT 174.520 56.450 175.865 56.680 ;
        RECT 176.370 56.540 178.940 57.360 ;
        RECT 179.120 56.680 181.860 57.360 ;
        RECT 181.880 56.550 183.710 57.360 ;
        RECT 184.635 57.130 186.325 57.360 ;
        RECT 176.370 56.450 177.960 56.540 ;
        RECT 184.635 56.450 186.470 57.130 ;
        RECT 186.480 56.550 187.850 57.360 ;
        RECT 187.870 56.490 188.300 57.275 ;
        RECT 188.320 56.680 191.990 57.360 ;
        RECT 188.320 56.450 189.250 56.680 ;
        RECT 192.000 56.580 193.370 57.360 ;
        RECT 194.300 56.680 203.490 57.360 ;
        RECT 198.810 56.460 199.740 56.680 ;
        RECT 202.570 56.450 203.490 56.680 ;
        RECT 203.810 56.680 205.645 57.360 ;
        RECT 203.810 56.450 204.740 56.680 ;
        RECT 205.800 56.550 208.550 57.360 ;
        RECT 209.330 56.680 211.165 57.360 ;
        RECT 211.465 57.360 211.630 57.380 ;
        RECT 214.220 57.360 214.390 57.550 ;
        RECT 217.450 57.405 217.610 57.515 ;
        RECT 222.315 57.380 222.485 57.570 ;
        RECT 227.100 57.520 227.270 57.550 ;
        RECT 226.175 57.410 226.295 57.520 ;
        RECT 227.095 57.410 227.270 57.520 ;
        RECT 227.100 57.360 227.270 57.410 ;
        RECT 227.560 57.360 227.730 57.570 ;
        RECT 231.240 57.380 231.410 57.570 ;
        RECT 236.760 57.380 236.930 57.550 ;
        RECT 239.055 57.410 239.175 57.520 ;
        RECT 240.440 57.380 240.610 57.570 ;
        RECT 242.280 57.380 242.450 57.570 ;
        RECT 236.765 57.360 236.930 57.380 ;
        RECT 243.200 57.360 243.370 57.550 ;
        RECT 245.500 57.380 245.670 57.550 ;
        RECT 245.500 57.360 245.665 57.380 ;
        RECT 245.960 57.360 246.130 57.570 ;
        RECT 247.340 57.360 247.510 57.550 ;
        RECT 251.490 57.415 251.650 57.525 ;
        RECT 252.860 57.380 253.030 57.570 ;
        RECT 253.780 57.360 253.950 57.550 ;
        RECT 254.240 57.360 254.410 57.550 ;
        RECT 263.440 57.360 263.610 57.550 ;
        RECT 264.820 57.520 264.990 57.570 ;
        RECT 264.815 57.410 264.990 57.520 ;
        RECT 264.820 57.380 264.990 57.410 ;
        RECT 265.280 57.380 265.450 57.570 ;
        RECT 265.740 57.360 265.910 57.550 ;
        RECT 268.960 57.380 269.130 57.570 ;
        RECT 274.480 57.550 274.620 57.570 ;
        RECT 271.260 57.360 271.430 57.550 ;
        RECT 274.480 57.380 274.650 57.550 ;
        RECT 274.940 57.520 275.110 57.570 ;
        RECT 274.935 57.410 275.110 57.520 ;
        RECT 274.940 57.380 275.110 57.410 ;
        RECT 275.400 57.360 275.570 57.550 ;
        RECT 277.695 57.410 277.815 57.520 ;
        RECT 278.895 57.380 279.065 57.570 ;
        RECT 282.755 57.410 282.875 57.520 ;
        RECT 283.220 57.380 283.390 57.570 ;
        RECT 289.200 57.360 289.370 57.550 ;
        RECT 289.660 57.360 289.830 57.550 ;
        RECT 291.775 57.360 291.945 57.550 ;
        RECT 292.880 57.380 293.050 57.570 ;
        RECT 295.640 57.360 295.810 57.550 ;
        RECT 299.315 57.410 299.435 57.520 ;
        RECT 303.460 57.380 303.630 57.570 ;
        RECT 304.380 57.380 304.550 57.570 ;
        RECT 308.980 57.360 309.150 57.550 ;
        RECT 309.435 57.410 309.555 57.520 ;
        RECT 310.820 57.360 310.990 57.570 ;
        RECT 211.465 56.680 213.300 57.360 ;
        RECT 209.330 56.450 210.260 56.680 ;
        RECT 212.370 56.450 213.300 56.680 ;
        RECT 213.630 56.490 214.060 57.275 ;
        RECT 214.160 56.450 217.160 57.360 ;
        RECT 218.220 56.680 227.410 57.360 ;
        RECT 227.420 56.680 236.610 57.360 ;
        RECT 236.765 56.680 238.600 57.360 ;
        RECT 218.220 56.450 219.140 56.680 ;
        RECT 221.970 56.460 222.900 56.680 ;
        RECT 231.930 56.460 232.860 56.680 ;
        RECT 235.690 56.450 236.610 56.680 ;
        RECT 237.670 56.450 238.600 56.680 ;
        RECT 239.390 56.490 239.820 57.275 ;
        RECT 239.935 56.680 243.400 57.360 ;
        RECT 243.830 56.680 245.665 57.360 ;
        RECT 239.935 56.450 240.855 56.680 ;
        RECT 243.830 56.450 244.760 56.680 ;
        RECT 245.820 56.550 247.190 57.360 ;
        RECT 247.310 56.680 250.775 57.360 ;
        RECT 249.855 56.450 250.775 56.680 ;
        RECT 250.880 56.450 254.090 57.360 ;
        RECT 254.100 56.680 263.290 57.360 ;
        RECT 258.610 56.460 259.540 56.680 ;
        RECT 262.370 56.450 263.290 56.680 ;
        RECT 263.310 56.450 264.660 57.360 ;
        RECT 265.150 56.490 265.580 57.275 ;
        RECT 265.600 56.550 271.110 57.360 ;
        RECT 271.120 56.550 274.790 57.360 ;
        RECT 275.260 56.680 284.450 57.360 ;
        RECT 284.695 56.680 289.510 57.360 ;
        RECT 279.770 56.460 280.700 56.680 ;
        RECT 283.530 56.450 284.450 56.680 ;
        RECT 289.520 56.550 290.890 57.360 ;
        RECT 290.910 56.490 291.340 57.275 ;
        RECT 291.360 56.680 295.260 57.360 ;
        RECT 291.360 56.450 292.290 56.680 ;
        RECT 295.500 56.550 299.170 57.360 ;
        RECT 299.645 56.680 309.290 57.360 ;
        RECT 299.645 56.560 302.345 56.680 ;
        RECT 299.645 56.450 301.415 56.560 ;
        RECT 307.010 56.460 307.930 56.680 ;
        RECT 309.760 56.550 311.130 57.360 ;
      LAYER nwell ;
        RECT 161.905 53.330 311.325 56.160 ;
      LAYER pwell ;
        RECT 162.100 52.130 163.470 52.940 ;
        RECT 163.480 52.130 165.310 52.940 ;
        RECT 170.290 52.810 171.220 53.030 ;
        RECT 174.050 52.810 174.970 53.040 ;
        RECT 165.780 52.130 174.970 52.810 ;
        RECT 174.990 52.215 175.420 53.000 ;
        RECT 175.440 52.810 176.370 53.040 ;
        RECT 184.875 52.810 186.010 53.040 ;
        RECT 175.440 52.130 179.340 52.810 ;
        RECT 179.590 52.130 182.330 52.810 ;
        RECT 182.800 52.130 186.010 52.810 ;
        RECT 186.020 52.840 186.950 53.040 ;
        RECT 188.280 52.840 189.230 53.040 ;
        RECT 186.020 52.360 189.230 52.840 ;
        RECT 186.165 52.160 189.230 52.360 ;
        RECT 162.240 51.920 162.410 52.130 ;
        RECT 163.620 51.920 163.790 52.130 ;
        RECT 165.455 51.970 165.575 52.080 ;
        RECT 165.920 51.920 166.090 52.130 ;
        RECT 175.120 51.920 175.290 52.110 ;
        RECT 175.855 51.940 176.025 52.130 ;
        RECT 182.020 51.940 182.190 52.130 ;
        RECT 182.475 51.970 182.595 52.080 ;
        RECT 182.940 51.940 183.110 52.130 ;
        RECT 186.165 51.940 186.335 52.160 ;
        RECT 188.295 52.130 189.230 52.160 ;
        RECT 189.990 52.130 192.910 53.040 ;
        RECT 193.155 52.130 197.970 52.810 ;
        RECT 197.980 52.130 200.170 53.040 ;
        RECT 200.750 52.215 201.180 53.000 ;
        RECT 201.200 52.130 202.570 52.940 ;
        RECT 202.890 52.810 203.820 53.040 ;
        RECT 206.020 52.950 206.970 53.040 ;
        RECT 202.890 52.130 204.725 52.810 ;
        RECT 187.540 51.920 187.710 52.110 ;
        RECT 189.380 52.080 189.550 52.110 ;
        RECT 188.470 51.965 188.630 52.075 ;
        RECT 189.375 51.970 189.550 52.080 ;
        RECT 189.380 51.920 189.550 51.970 ;
        RECT 192.595 52.075 192.765 52.130 ;
        RECT 192.595 51.965 192.770 52.075 ;
        RECT 192.595 51.940 192.765 51.965 ;
        RECT 193.520 51.940 193.690 52.110 ;
        RECT 195.360 51.920 195.530 52.110 ;
        RECT 197.660 51.940 197.830 52.130 ;
        RECT 198.125 51.940 198.295 52.130 ;
        RECT 200.415 51.970 200.535 52.080 ;
        RECT 201.340 51.940 201.510 52.130 ;
        RECT 204.560 52.110 204.725 52.130 ;
        RECT 205.040 52.130 206.970 52.950 ;
        RECT 207.180 52.130 209.930 52.940 ;
        RECT 214.450 52.810 215.380 53.030 ;
        RECT 218.210 52.810 219.130 53.040 ;
        RECT 220.190 52.810 221.120 53.040 ;
        RECT 209.940 52.130 219.130 52.810 ;
        RECT 219.285 52.130 221.120 52.810 ;
        RECT 221.440 52.130 226.255 52.810 ;
        RECT 226.510 52.215 226.940 53.000 ;
        RECT 226.960 52.130 237.970 53.040 ;
        RECT 238.325 52.130 241.980 53.040 ;
        RECT 242.235 52.810 243.155 53.040 ;
        RECT 248.475 52.810 249.395 53.040 ;
        RECT 242.235 52.130 245.700 52.810 ;
        RECT 245.930 52.130 249.395 52.810 ;
        RECT 249.500 52.130 252.250 52.940 ;
        RECT 252.270 52.215 252.700 53.000 ;
        RECT 263.855 52.810 264.775 53.040 ;
        RECT 253.875 52.130 258.690 52.810 ;
        RECT 258.935 52.130 263.750 52.810 ;
        RECT 263.855 52.130 267.320 52.810 ;
        RECT 267.440 52.130 271.095 53.040 ;
        RECT 271.120 52.130 274.790 52.940 ;
        RECT 274.850 52.130 278.010 53.040 ;
        RECT 278.030 52.215 278.460 53.000 ;
        RECT 278.480 52.810 279.400 53.040 ;
        RECT 282.230 52.810 283.160 53.030 ;
        RECT 278.480 52.130 287.670 52.810 ;
        RECT 287.680 52.130 292.495 52.810 ;
        RECT 292.740 52.130 298.250 52.940 ;
        RECT 298.260 52.130 301.010 52.940 ;
        RECT 301.020 52.130 303.760 52.810 ;
        RECT 303.790 52.215 304.220 53.000 ;
        RECT 306.895 52.810 307.815 53.040 ;
        RECT 304.350 52.130 307.815 52.810 ;
        RECT 308.380 52.130 309.750 52.910 ;
        RECT 309.760 52.130 311.130 52.940 ;
        RECT 205.040 52.110 205.190 52.130 ;
        RECT 204.560 51.920 204.730 52.110 ;
        RECT 205.020 51.940 205.190 52.110 ;
        RECT 207.320 51.940 207.490 52.130 ;
        RECT 210.080 51.940 210.250 52.130 ;
        RECT 219.285 52.110 219.450 52.130 ;
        RECT 214.220 51.920 214.390 52.110 ;
        RECT 219.280 51.940 219.450 52.110 ;
        RECT 221.580 51.940 221.750 52.130 ;
        RECT 223.420 51.920 223.590 52.110 ;
        RECT 227.105 51.940 227.275 52.130 ;
        RECT 241.820 52.110 241.980 52.130 ;
        RECT 228.480 51.920 228.650 52.110 ;
        RECT 230.320 51.920 230.490 52.110 ;
        RECT 241.820 51.940 241.990 52.110 ;
        RECT 243.660 51.940 243.830 52.110 ;
        RECT 243.660 51.920 243.820 51.940 ;
        RECT 244.120 51.920 244.290 52.110 ;
        RECT 245.500 51.940 245.670 52.130 ;
        RECT 245.960 51.940 246.130 52.130 ;
        RECT 249.640 51.940 249.810 52.130 ;
        RECT 250.560 51.940 250.730 52.110 ;
        RECT 252.870 51.975 253.030 52.085 ;
        RECT 250.560 51.920 250.720 51.940 ;
        RECT 254.240 51.920 254.410 52.110 ;
        RECT 254.700 51.920 254.870 52.110 ;
        RECT 256.080 51.920 256.250 52.110 ;
        RECT 258.380 51.940 258.550 52.130 ;
        RECT 263.440 51.940 263.610 52.130 ;
        RECT 265.740 51.920 265.910 52.110 ;
        RECT 267.120 51.940 267.290 52.130 ;
        RECT 267.585 52.080 267.755 52.130 ;
        RECT 267.575 51.970 267.755 52.080 ;
        RECT 267.585 51.940 267.755 51.970 ;
        RECT 268.040 51.920 268.210 52.110 ;
        RECT 271.260 51.940 271.430 52.130 ;
        RECT 274.940 51.940 275.110 52.130 ;
        RECT 285.980 51.920 286.150 52.110 ;
        RECT 287.360 51.940 287.530 52.130 ;
        RECT 287.820 51.940 287.990 52.130 ;
        RECT 289.660 51.920 289.830 52.110 ;
        RECT 290.130 51.965 290.290 52.075 ;
        RECT 291.500 51.940 291.670 52.110 ;
        RECT 292.880 51.940 293.050 52.130 ;
        RECT 294.720 51.920 294.890 52.110 ;
        RECT 298.400 51.920 298.570 52.130 ;
        RECT 301.160 51.940 301.330 52.130 ;
        RECT 304.380 51.940 304.550 52.130 ;
        RECT 308.055 51.970 308.175 52.080 ;
        RECT 308.980 51.920 309.150 52.110 ;
        RECT 309.440 52.080 309.610 52.130 ;
        RECT 309.435 51.970 309.610 52.080 ;
        RECT 309.440 51.940 309.610 51.970 ;
        RECT 310.820 51.920 310.990 52.130 ;
        RECT 162.100 51.110 163.470 51.920 ;
        RECT 163.480 51.110 165.310 51.920 ;
        RECT 165.780 51.240 174.970 51.920 ;
        RECT 174.980 51.240 184.170 51.920 ;
        RECT 170.290 51.020 171.220 51.240 ;
        RECT 174.050 51.010 174.970 51.240 ;
        RECT 179.490 51.020 180.420 51.240 ;
        RECT 183.250 51.010 184.170 51.240 ;
        RECT 184.180 51.240 187.850 51.920 ;
        RECT 184.180 51.010 185.110 51.240 ;
        RECT 187.870 51.050 188.300 51.835 ;
        RECT 189.240 51.240 192.450 51.920 ;
        RECT 193.845 51.240 195.210 51.920 ;
        RECT 195.220 51.240 204.410 51.920 ;
        RECT 204.420 51.240 213.610 51.920 ;
        RECT 191.315 51.010 192.450 51.240 ;
        RECT 199.730 51.020 200.660 51.240 ;
        RECT 203.490 51.010 204.410 51.240 ;
        RECT 208.930 51.020 209.860 51.240 ;
        RECT 212.690 51.010 213.610 51.240 ;
        RECT 213.630 51.050 214.060 51.835 ;
        RECT 214.080 51.240 223.270 51.920 ;
        RECT 223.280 51.240 228.095 51.920 ;
        RECT 218.590 51.020 219.520 51.240 ;
        RECT 222.350 51.010 223.270 51.240 ;
        RECT 228.340 51.110 230.170 51.920 ;
        RECT 230.180 51.240 239.370 51.920 ;
        RECT 234.690 51.020 235.620 51.240 ;
        RECT 238.450 51.010 239.370 51.240 ;
        RECT 239.390 51.050 239.820 51.835 ;
        RECT 240.165 51.010 243.820 51.920 ;
        RECT 243.980 51.110 246.730 51.920 ;
        RECT 247.065 51.010 250.720 51.920 ;
        RECT 250.975 51.240 254.440 51.920 ;
        RECT 250.975 51.010 251.895 51.240 ;
        RECT 254.560 51.110 255.930 51.920 ;
        RECT 255.940 51.240 265.130 51.920 ;
        RECT 260.450 51.020 261.380 51.240 ;
        RECT 264.210 51.010 265.130 51.240 ;
        RECT 265.150 51.050 265.580 51.835 ;
        RECT 265.600 51.110 267.430 51.920 ;
        RECT 267.900 51.240 277.090 51.920 ;
        RECT 272.410 51.020 273.340 51.240 ;
        RECT 276.170 51.010 277.090 51.240 ;
        RECT 277.100 51.240 286.290 51.920 ;
        RECT 286.395 51.240 289.860 51.920 ;
        RECT 277.100 51.010 278.020 51.240 ;
        RECT 280.850 51.020 281.780 51.240 ;
        RECT 286.395 51.010 287.315 51.240 ;
        RECT 290.910 51.050 291.340 51.835 ;
        RECT 291.765 51.240 294.190 51.920 ;
        RECT 294.580 51.110 298.250 51.920 ;
        RECT 298.260 51.110 299.630 51.920 ;
        RECT 300.010 51.240 309.290 51.920 ;
        RECT 300.010 51.120 302.345 51.240 ;
        RECT 300.010 51.010 300.930 51.120 ;
        RECT 307.010 51.020 307.930 51.240 ;
        RECT 309.760 51.110 311.130 51.920 ;
      LAYER nwell ;
        RECT 161.905 47.890 311.325 50.720 ;
      LAYER pwell ;
        RECT 162.100 46.690 163.470 47.500 ;
        RECT 163.480 46.690 168.990 47.500 ;
        RECT 169.000 46.690 174.510 47.500 ;
        RECT 174.990 46.775 175.420 47.560 ;
        RECT 175.440 47.370 176.370 47.600 ;
        RECT 179.580 47.370 180.510 47.600 ;
        RECT 175.440 46.690 179.340 47.370 ;
        RECT 179.580 46.690 183.480 47.370 ;
        RECT 184.200 46.690 185.550 47.600 ;
        RECT 185.560 46.690 188.310 47.500 ;
        RECT 188.330 46.690 189.680 47.600 ;
        RECT 189.700 46.690 193.370 47.500 ;
        RECT 193.380 46.690 194.750 47.500 ;
        RECT 194.995 46.690 199.810 47.370 ;
        RECT 200.750 46.775 201.180 47.560 ;
        RECT 201.200 46.690 206.710 47.500 ;
        RECT 206.720 46.690 212.230 47.500 ;
        RECT 212.240 46.690 214.070 47.500 ;
        RECT 214.390 47.370 215.320 47.600 ;
        RECT 220.890 47.370 221.820 47.590 ;
        RECT 224.650 47.370 225.570 47.600 ;
        RECT 214.390 46.690 216.225 47.370 ;
        RECT 216.380 46.690 225.570 47.370 ;
        RECT 226.510 46.775 226.940 47.560 ;
        RECT 226.960 46.690 228.330 47.500 ;
        RECT 230.995 47.370 231.915 47.600 ;
        RECT 236.530 47.370 237.460 47.590 ;
        RECT 240.290 47.370 241.210 47.600 ;
        RECT 228.450 46.690 231.915 47.370 ;
        RECT 232.020 46.690 241.210 47.370 ;
        RECT 241.220 47.370 242.140 47.600 ;
        RECT 244.970 47.370 245.900 47.590 ;
        RECT 241.220 46.690 250.410 47.370 ;
        RECT 250.420 46.690 252.250 47.500 ;
        RECT 252.270 46.775 252.700 47.560 ;
        RECT 252.770 46.690 255.930 47.600 ;
        RECT 260.450 47.370 261.380 47.590 ;
        RECT 264.210 47.370 265.130 47.600 ;
        RECT 266.510 47.370 267.430 47.600 ;
        RECT 255.940 46.690 265.130 47.370 ;
        RECT 265.140 46.690 267.430 47.370 ;
        RECT 267.455 47.370 268.825 47.600 ;
        RECT 267.455 46.690 269.730 47.370 ;
        RECT 269.840 46.690 272.030 47.600 ;
        RECT 272.040 46.690 277.550 47.500 ;
        RECT 278.030 46.775 278.460 47.560 ;
        RECT 281.680 47.370 282.610 47.600 ;
        RECT 288.050 47.370 288.980 47.590 ;
        RECT 291.810 47.370 292.730 47.600 ;
        RECT 278.710 46.690 282.610 47.370 ;
        RECT 283.540 46.690 292.730 47.370 ;
        RECT 292.835 47.370 293.755 47.600 ;
        RECT 292.835 46.690 296.300 47.370 ;
        RECT 296.420 46.690 301.930 47.500 ;
        RECT 301.940 46.690 303.770 47.500 ;
        RECT 303.790 46.775 304.220 47.560 ;
        RECT 304.240 46.690 309.750 47.500 ;
        RECT 309.760 46.690 311.130 47.500 ;
        RECT 162.240 46.480 162.410 46.690 ;
        RECT 163.620 46.480 163.790 46.690 ;
        RECT 169.140 46.480 169.310 46.690 ;
        RECT 172.820 46.480 172.990 46.670 ;
        RECT 174.655 46.530 174.775 46.640 ;
        RECT 175.855 46.500 176.025 46.690 ;
        RECT 179.995 46.500 180.165 46.690 ;
        RECT 183.855 46.530 183.975 46.640 ;
        RECT 185.235 46.500 185.405 46.690 ;
        RECT 185.700 46.480 185.870 46.690 ;
        RECT 186.160 46.480 186.330 46.670 ;
        RECT 188.460 46.500 188.630 46.690 ;
        RECT 189.840 46.480 190.010 46.690 ;
        RECT 190.300 46.480 190.470 46.670 ;
        RECT 193.520 46.500 193.690 46.690 ;
        RECT 199.500 46.500 199.670 46.690 ;
        RECT 199.970 46.525 200.130 46.645 ;
        RECT 200.885 46.480 201.055 46.670 ;
        RECT 201.340 46.500 201.510 46.690 ;
        RECT 204.100 46.480 204.270 46.670 ;
        RECT 206.860 46.500 207.030 46.690 ;
        RECT 209.620 46.480 209.790 46.670 ;
        RECT 212.380 46.500 212.550 46.690 ;
        RECT 216.060 46.670 216.225 46.690 ;
        RECT 213.295 46.530 213.415 46.640 ;
        RECT 214.220 46.480 214.390 46.670 ;
        RECT 216.060 46.640 216.230 46.670 ;
        RECT 216.055 46.530 216.230 46.640 ;
        RECT 216.060 46.500 216.230 46.530 ;
        RECT 216.520 46.500 216.690 46.690 ;
        RECT 216.795 46.480 216.965 46.670 ;
        RECT 220.670 46.525 220.830 46.635 ;
        RECT 224.340 46.500 224.510 46.670 ;
        RECT 225.730 46.535 225.890 46.645 ;
        RECT 227.100 46.500 227.270 46.690 ;
        RECT 228.020 46.480 228.190 46.670 ;
        RECT 228.480 46.480 228.650 46.690 ;
        RECT 230.320 46.480 230.490 46.670 ;
        RECT 232.160 46.500 232.330 46.690 ;
        RECT 243.660 46.500 243.830 46.670 ;
        RECT 243.660 46.480 243.820 46.500 ;
        RECT 247.340 46.480 247.510 46.670 ;
        RECT 247.795 46.530 247.915 46.640 ;
        RECT 248.260 46.480 248.430 46.670 ;
        RECT 250.100 46.500 250.270 46.690 ;
        RECT 250.560 46.500 250.730 46.690 ;
        RECT 252.860 46.500 253.030 46.690 ;
        RECT 256.080 46.500 256.250 46.690 ;
        RECT 261.140 46.500 261.310 46.670 ;
        RECT 261.140 46.480 261.300 46.500 ;
        RECT 264.820 46.480 264.990 46.670 ;
        RECT 265.280 46.500 265.450 46.690 ;
        RECT 269.415 46.670 269.585 46.690 ;
        RECT 271.715 46.670 271.885 46.690 ;
        RECT 267.580 46.500 267.750 46.670 ;
        RECT 267.580 46.480 267.745 46.500 ;
        RECT 268.040 46.480 268.210 46.670 ;
        RECT 269.415 46.500 269.590 46.670 ;
        RECT 271.255 46.530 271.375 46.640 ;
        RECT 271.715 46.500 271.895 46.670 ;
        RECT 272.180 46.500 272.350 46.690 ;
        RECT 273.555 46.530 273.675 46.640 ;
        RECT 269.420 46.480 269.590 46.500 ;
        RECT 271.725 46.480 271.895 46.500 ;
        RECT 277.240 46.480 277.410 46.670 ;
        RECT 277.700 46.640 277.870 46.670 ;
        RECT 277.695 46.530 277.870 46.640 ;
        RECT 277.700 46.480 277.870 46.530 ;
        RECT 279.080 46.480 279.250 46.670 ;
        RECT 282.025 46.500 282.195 46.690 ;
        RECT 282.760 46.480 282.930 46.670 ;
        RECT 283.680 46.500 283.850 46.690 ;
        RECT 288.280 46.480 288.450 46.670 ;
        RECT 291.500 46.480 291.670 46.670 ;
        RECT 295.180 46.480 295.350 46.670 ;
        RECT 296.100 46.500 296.270 46.690 ;
        RECT 296.560 46.480 296.730 46.690 ;
        RECT 302.080 46.500 302.250 46.690 ;
        RECT 304.380 46.500 304.550 46.690 ;
        RECT 305.760 46.480 305.930 46.670 ;
        RECT 307.595 46.530 307.715 46.640 ;
        RECT 308.060 46.480 308.230 46.670 ;
        RECT 310.820 46.480 310.990 46.690 ;
        RECT 162.100 45.670 163.470 46.480 ;
        RECT 163.480 45.670 168.990 46.480 ;
        RECT 169.000 45.670 172.670 46.480 ;
        RECT 172.680 45.800 182.290 46.480 ;
        RECT 177.190 45.580 178.120 45.800 ;
        RECT 180.950 45.570 182.290 45.800 ;
        RECT 182.435 45.800 185.900 46.480 ;
        RECT 182.435 45.570 183.355 45.800 ;
        RECT 186.020 45.670 187.850 46.480 ;
        RECT 187.870 45.610 188.300 46.395 ;
        RECT 188.320 45.800 190.150 46.480 ;
        RECT 190.160 45.800 199.770 46.480 ;
        RECT 200.740 45.800 203.950 46.480 ;
        RECT 194.670 45.580 195.600 45.800 ;
        RECT 198.430 45.570 199.770 45.800 ;
        RECT 202.585 45.570 203.950 45.800 ;
        RECT 203.960 45.670 209.470 46.480 ;
        RECT 209.480 45.670 213.150 46.480 ;
        RECT 213.630 45.610 214.060 46.395 ;
        RECT 214.080 45.670 215.910 46.480 ;
        RECT 216.380 45.800 220.280 46.480 ;
        RECT 221.820 45.800 224.245 46.480 ;
        RECT 224.755 45.800 228.220 46.480 ;
        RECT 228.340 45.800 230.170 46.480 ;
        RECT 230.180 45.800 239.370 46.480 ;
        RECT 216.380 45.570 217.310 45.800 ;
        RECT 224.755 45.570 225.675 45.800 ;
        RECT 228.825 45.570 230.170 45.800 ;
        RECT 234.690 45.580 235.620 45.800 ;
        RECT 238.450 45.570 239.370 45.800 ;
        RECT 239.390 45.610 239.820 46.395 ;
        RECT 240.165 45.570 243.820 46.480 ;
        RECT 244.075 45.800 247.540 46.480 ;
        RECT 248.120 45.800 257.310 46.480 ;
        RECT 244.075 45.570 244.995 45.800 ;
        RECT 252.630 45.580 253.560 45.800 ;
        RECT 256.390 45.570 257.310 45.800 ;
        RECT 257.645 45.570 261.300 46.480 ;
        RECT 261.555 45.800 265.020 46.480 ;
        RECT 261.555 45.570 262.475 45.800 ;
        RECT 265.150 45.610 265.580 46.395 ;
        RECT 265.910 45.800 267.745 46.480 ;
        RECT 265.910 45.570 266.840 45.800 ;
        RECT 267.910 45.570 269.260 46.480 ;
        RECT 269.280 45.670 271.110 46.480 ;
        RECT 271.580 45.570 273.410 46.480 ;
        RECT 273.975 45.800 277.440 46.480 ;
        RECT 273.975 45.570 274.895 45.800 ;
        RECT 277.560 45.670 278.930 46.480 ;
        RECT 279.050 45.800 282.515 46.480 ;
        RECT 281.595 45.570 282.515 45.800 ;
        RECT 282.620 45.670 288.130 46.480 ;
        RECT 288.140 45.670 290.890 46.480 ;
        RECT 290.910 45.610 291.340 46.395 ;
        RECT 291.360 45.670 295.030 46.480 ;
        RECT 295.040 45.670 296.410 46.480 ;
        RECT 296.420 45.800 305.610 46.480 ;
        RECT 300.930 45.580 301.860 45.800 ;
        RECT 304.690 45.570 305.610 45.800 ;
        RECT 305.620 45.670 307.450 46.480 ;
        RECT 307.920 45.800 309.750 46.480 ;
        RECT 308.405 45.570 309.750 45.800 ;
        RECT 309.760 45.670 311.130 46.480 ;
      LAYER nwell ;
        RECT 161.905 42.450 311.325 45.280 ;
      LAYER pwell ;
        RECT 162.100 41.250 163.470 42.060 ;
        RECT 163.480 41.250 165.310 42.060 ;
        RECT 170.290 41.930 171.220 42.150 ;
        RECT 174.050 41.930 174.970 42.160 ;
        RECT 165.780 41.250 174.970 41.930 ;
        RECT 174.990 41.335 175.420 42.120 ;
        RECT 179.950 41.930 180.880 42.150 ;
        RECT 183.710 41.930 184.630 42.160 ;
        RECT 175.440 41.250 184.630 41.930 ;
        RECT 184.640 41.250 186.470 42.060 ;
        RECT 186.520 41.930 187.860 42.160 ;
        RECT 190.690 41.930 191.620 42.150 ;
        RECT 186.520 41.250 196.130 41.930 ;
        RECT 196.140 41.250 199.810 42.060 ;
        RECT 200.750 41.335 201.180 42.120 ;
        RECT 205.710 41.930 206.640 42.150 ;
        RECT 209.470 41.930 210.390 42.160 ;
        RECT 201.200 41.250 210.390 41.930 ;
        RECT 210.495 41.930 211.415 42.160 ;
        RECT 219.510 41.930 220.440 42.150 ;
        RECT 223.270 41.930 224.610 42.160 ;
        RECT 210.495 41.250 213.960 41.930 ;
        RECT 215.000 41.250 224.610 41.930 ;
        RECT 224.660 41.250 226.490 42.060 ;
        RECT 226.510 41.335 226.940 42.120 ;
        RECT 230.735 41.930 231.655 42.160 ;
        RECT 226.970 41.250 229.710 41.930 ;
        RECT 230.735 41.250 234.200 41.930 ;
        RECT 235.105 41.250 238.760 42.160 ;
        RECT 238.920 41.250 240.290 42.060 ;
        RECT 240.300 41.930 241.230 42.160 ;
        RECT 247.095 41.930 248.015 42.160 ;
        RECT 240.300 41.250 244.200 41.930 ;
        RECT 244.550 41.250 248.015 41.930 ;
        RECT 248.430 41.930 249.360 42.160 ;
        RECT 248.430 41.250 250.265 41.930 ;
        RECT 250.420 41.250 252.250 42.060 ;
        RECT 252.270 41.335 252.700 42.120 ;
        RECT 256.250 41.930 257.180 42.160 ;
        RECT 253.125 41.250 255.550 41.930 ;
        RECT 256.250 41.250 258.085 41.930 ;
        RECT 259.180 41.250 260.530 42.160 ;
        RECT 260.540 41.250 264.210 42.060 ;
        RECT 264.220 41.250 265.590 42.060 ;
        RECT 270.110 41.930 271.040 42.150 ;
        RECT 273.870 41.930 274.790 42.160 ;
        RECT 265.600 41.250 274.790 41.930 ;
        RECT 274.810 41.250 277.550 41.930 ;
        RECT 278.030 41.335 278.460 42.120 ;
        RECT 278.575 41.930 279.495 42.160 ;
        RECT 278.575 41.250 282.040 41.930 ;
        RECT 282.160 41.250 284.910 42.060 ;
        RECT 285.380 41.930 286.300 42.160 ;
        RECT 289.130 41.930 290.060 42.150 ;
        RECT 285.380 41.250 294.570 41.930 ;
        RECT 294.580 41.250 300.090 42.060 ;
        RECT 300.100 41.250 303.770 42.060 ;
        RECT 303.790 41.335 304.220 42.120 ;
        RECT 308.735 41.930 309.655 42.160 ;
        RECT 304.240 41.250 306.070 41.930 ;
        RECT 306.190 41.250 309.655 41.930 ;
        RECT 309.760 41.250 311.130 42.060 ;
        RECT 162.240 41.040 162.410 41.250 ;
        RECT 163.620 41.040 163.790 41.250 ;
        RECT 165.455 41.090 165.575 41.200 ;
        RECT 165.920 41.060 166.090 41.250 ;
        RECT 167.310 41.085 167.470 41.195 ;
        RECT 168.220 41.040 168.390 41.230 ;
        RECT 175.580 41.060 175.750 41.250 ;
        RECT 177.695 41.040 177.865 41.230 ;
        RECT 181.560 41.040 181.730 41.230 ;
        RECT 183.395 41.090 183.515 41.200 ;
        RECT 184.135 41.040 184.305 41.230 ;
        RECT 184.780 41.060 184.950 41.250 ;
        RECT 188.460 41.040 188.630 41.230 ;
        RECT 190.115 41.040 190.285 41.230 ;
        RECT 193.980 41.040 194.150 41.230 ;
        RECT 195.360 41.040 195.530 41.230 ;
        RECT 195.820 41.060 195.990 41.250 ;
        RECT 196.280 41.060 196.450 41.250 ;
        RECT 199.970 41.095 200.130 41.205 ;
        RECT 201.340 41.060 201.510 41.250 ;
        RECT 204.835 41.040 205.005 41.230 ;
        RECT 208.700 41.040 208.870 41.230 ;
        RECT 210.080 41.040 210.250 41.230 ;
        RECT 213.760 41.060 213.930 41.250 ;
        RECT 214.220 41.040 214.390 41.230 ;
        RECT 215.140 41.060 215.310 41.250 ;
        RECT 224.800 41.060 224.970 41.250 ;
        RECT 225.260 41.060 225.430 41.230 ;
        RECT 225.260 41.040 225.425 41.060 ;
        RECT 225.995 41.040 226.165 41.230 ;
        RECT 229.400 41.060 229.570 41.250 ;
        RECT 229.870 41.095 230.030 41.205 ;
        RECT 230.135 41.040 230.305 41.230 ;
        RECT 234.000 41.040 234.170 41.250 ;
        RECT 238.600 41.230 238.760 41.250 ;
        RECT 234.455 41.090 234.575 41.200 ;
        RECT 238.600 41.060 238.770 41.230 ;
        RECT 239.060 41.040 239.230 41.250 ;
        RECT 239.980 41.040 240.150 41.230 ;
        RECT 240.715 41.060 240.885 41.250 ;
        RECT 241.635 41.040 241.805 41.230 ;
        RECT 244.580 41.060 244.750 41.250 ;
        RECT 250.100 41.230 250.265 41.250 ;
        RECT 245.775 41.040 245.945 41.230 ;
        RECT 250.100 41.060 250.270 41.230 ;
        RECT 250.560 41.060 250.730 41.250 ;
        RECT 257.920 41.230 258.085 41.250 ;
        RECT 252.860 41.040 253.030 41.230 ;
        RECT 253.320 41.040 253.490 41.230 ;
        RECT 254.700 41.040 254.870 41.230 ;
        RECT 257.920 41.060 258.090 41.230 ;
        RECT 258.390 41.095 258.550 41.205 ;
        RECT 259.295 41.060 259.465 41.250 ;
        RECT 260.680 41.230 260.850 41.250 ;
        RECT 260.675 41.060 260.850 41.230 ;
        RECT 260.675 41.040 260.845 41.060 ;
        RECT 261.140 41.040 261.310 41.230 ;
        RECT 263.900 41.040 264.070 41.230 ;
        RECT 264.360 41.060 264.530 41.250 ;
        RECT 265.740 41.060 265.910 41.250 ;
        RECT 277.240 41.230 277.410 41.250 ;
        RECT 268.960 41.040 269.130 41.230 ;
        RECT 269.430 41.085 269.590 41.195 ;
        RECT 271.260 41.040 271.430 41.230 ;
        RECT 271.725 41.040 271.895 41.230 ;
        RECT 277.235 41.060 277.410 41.230 ;
        RECT 277.695 41.090 277.815 41.200 ;
        RECT 277.235 41.040 277.405 41.060 ;
        RECT 279.080 41.040 279.250 41.230 ;
        RECT 279.535 41.090 279.655 41.200 ;
        RECT 281.840 41.060 282.010 41.250 ;
        RECT 282.300 41.060 282.470 41.250 ;
        RECT 283.220 41.040 283.390 41.230 ;
        RECT 283.680 41.040 283.850 41.230 ;
        RECT 285.055 41.090 285.175 41.200 ;
        RECT 289.200 41.040 289.370 41.230 ;
        RECT 291.500 41.040 291.670 41.230 ;
        RECT 294.260 41.060 294.430 41.250 ;
        RECT 294.720 41.060 294.890 41.250 ;
        RECT 297.020 41.040 297.190 41.230 ;
        RECT 300.240 41.060 300.410 41.250 ;
        RECT 304.380 41.060 304.550 41.250 ;
        RECT 306.220 41.060 306.390 41.250 ;
        RECT 308.520 41.040 308.690 41.230 ;
        RECT 308.990 41.085 309.150 41.195 ;
        RECT 310.820 41.040 310.990 41.250 ;
        RECT 162.100 40.230 163.470 41.040 ;
        RECT 163.480 40.230 167.150 41.040 ;
        RECT 168.080 40.360 177.270 41.040 ;
        RECT 172.590 40.140 173.520 40.360 ;
        RECT 176.350 40.130 177.270 40.360 ;
        RECT 177.280 40.360 181.180 41.040 ;
        RECT 177.280 40.130 178.210 40.360 ;
        RECT 181.420 40.230 183.250 41.040 ;
        RECT 183.720 40.360 187.620 41.040 ;
        RECT 183.720 40.130 184.650 40.360 ;
        RECT 187.870 40.170 188.300 40.955 ;
        RECT 188.320 40.230 189.690 41.040 ;
        RECT 189.700 40.360 193.600 41.040 ;
        RECT 189.700 40.130 190.630 40.360 ;
        RECT 193.840 40.230 195.210 41.040 ;
        RECT 195.220 40.360 204.410 41.040 ;
        RECT 199.730 40.140 200.660 40.360 ;
        RECT 203.490 40.130 204.410 40.360 ;
        RECT 204.420 40.360 208.320 41.040 ;
        RECT 204.420 40.130 205.350 40.360 ;
        RECT 208.560 40.230 209.930 41.040 ;
        RECT 210.050 40.360 213.515 41.040 ;
        RECT 212.595 40.130 213.515 40.360 ;
        RECT 213.630 40.170 214.060 40.955 ;
        RECT 214.080 40.360 223.270 41.040 ;
        RECT 218.590 40.140 219.520 40.360 ;
        RECT 222.350 40.130 223.270 40.360 ;
        RECT 223.590 40.360 225.425 41.040 ;
        RECT 225.580 40.360 229.480 41.040 ;
        RECT 229.720 40.360 233.620 41.040 ;
        RECT 233.970 40.360 237.435 41.040 ;
        RECT 237.540 40.360 239.370 41.040 ;
        RECT 223.590 40.130 224.520 40.360 ;
        RECT 225.580 40.130 226.510 40.360 ;
        RECT 229.720 40.130 230.650 40.360 ;
        RECT 236.515 40.130 237.435 40.360 ;
        RECT 239.390 40.170 239.820 40.955 ;
        RECT 239.840 40.230 241.210 41.040 ;
        RECT 241.220 40.360 245.120 41.040 ;
        RECT 245.360 40.360 249.260 41.040 ;
        RECT 249.595 40.360 253.060 41.040 ;
        RECT 241.220 40.130 242.150 40.360 ;
        RECT 245.360 40.130 246.290 40.360 ;
        RECT 249.595 40.130 250.515 40.360 ;
        RECT 253.180 40.230 254.550 41.040 ;
        RECT 254.560 40.360 256.850 41.040 ;
        RECT 255.930 40.130 256.850 40.360 ;
        RECT 257.100 40.130 260.990 41.040 ;
        RECT 261.000 40.130 263.750 41.040 ;
        RECT 263.760 40.230 265.130 41.040 ;
        RECT 265.150 40.170 265.580 40.955 ;
        RECT 265.695 40.360 269.160 41.040 ;
        RECT 265.695 40.130 266.615 40.360 ;
        RECT 270.210 40.130 271.560 41.040 ;
        RECT 271.580 40.360 275.575 41.040 ;
        RECT 272.065 40.130 275.575 40.360 ;
        RECT 275.780 40.130 277.550 41.040 ;
        RECT 277.560 40.130 279.375 41.040 ;
        RECT 279.955 40.360 283.420 41.040 ;
        RECT 279.955 40.130 280.875 40.360 ;
        RECT 283.540 40.230 289.050 41.040 ;
        RECT 289.060 40.230 290.890 41.040 ;
        RECT 290.910 40.170 291.340 40.955 ;
        RECT 291.360 40.230 296.870 41.040 ;
        RECT 296.880 40.230 299.630 41.040 ;
        RECT 299.640 40.360 308.830 41.040 ;
        RECT 299.640 40.130 300.560 40.360 ;
        RECT 303.390 40.140 304.320 40.360 ;
        RECT 309.760 40.230 311.130 41.040 ;
      LAYER nwell ;
        RECT 161.905 37.010 311.325 39.840 ;
      LAYER pwell ;
        RECT 162.100 35.810 163.470 36.620 ;
        RECT 163.480 35.810 167.150 36.620 ;
        RECT 167.255 36.490 168.175 36.720 ;
        RECT 170.840 36.490 171.770 36.720 ;
        RECT 167.255 35.810 170.720 36.490 ;
        RECT 170.840 35.810 174.740 36.490 ;
        RECT 174.990 35.895 175.420 36.680 ;
        RECT 175.440 36.490 176.370 36.720 ;
        RECT 183.155 36.490 184.075 36.720 ;
        RECT 188.690 36.490 189.620 36.710 ;
        RECT 192.450 36.490 193.370 36.720 ;
        RECT 175.440 35.810 179.340 36.490 ;
        RECT 180.610 35.810 184.075 36.490 ;
        RECT 184.180 35.810 193.370 36.490 ;
        RECT 193.475 36.490 194.395 36.720 ;
        RECT 199.715 36.490 200.635 36.720 ;
        RECT 193.475 35.810 196.940 36.490 ;
        RECT 197.170 35.810 200.635 36.490 ;
        RECT 200.750 35.895 201.180 36.680 ;
        RECT 201.200 35.810 203.950 36.620 ;
        RECT 204.420 36.490 205.350 36.720 ;
        RECT 204.420 35.810 208.320 36.490 ;
        RECT 208.560 35.810 210.390 36.620 ;
        RECT 214.060 36.490 214.990 36.720 ;
        RECT 211.090 35.810 214.990 36.490 ;
        RECT 215.000 36.490 215.930 36.720 ;
        RECT 219.235 36.490 220.155 36.720 ;
        RECT 222.915 36.490 223.835 36.720 ;
        RECT 215.000 35.810 218.900 36.490 ;
        RECT 219.235 35.810 222.700 36.490 ;
        RECT 222.915 35.810 226.380 36.490 ;
        RECT 226.510 35.895 226.940 36.680 ;
        RECT 226.960 35.810 228.790 36.620 ;
        RECT 233.310 36.490 234.240 36.710 ;
        RECT 237.070 36.490 238.410 36.720 ;
        RECT 228.800 35.810 238.410 36.490 ;
        RECT 238.460 35.810 239.830 36.620 ;
        RECT 244.350 36.490 245.280 36.710 ;
        RECT 248.110 36.490 249.030 36.720 ;
        RECT 239.840 35.810 249.030 36.490 ;
        RECT 249.040 35.810 251.790 36.620 ;
        RECT 252.270 35.895 252.700 36.680 ;
        RECT 252.720 35.810 254.090 36.620 ;
        RECT 258.610 36.490 259.540 36.710 ;
        RECT 262.370 36.490 263.290 36.720 ;
        RECT 254.100 35.810 263.290 36.490 ;
        RECT 263.610 36.490 264.540 36.720 ;
        RECT 265.800 36.630 266.750 36.720 ;
        RECT 263.610 35.810 265.445 36.490 ;
        RECT 265.800 35.810 267.730 36.630 ;
        RECT 273.330 36.490 274.260 36.710 ;
        RECT 277.090 36.490 278.010 36.720 ;
        RECT 268.820 35.810 278.010 36.490 ;
        RECT 278.030 35.895 278.460 36.680 ;
        RECT 278.480 36.520 279.410 36.720 ;
        RECT 280.740 36.520 281.690 36.720 ;
        RECT 278.480 36.040 281.690 36.520 ;
        RECT 278.625 35.840 281.690 36.040 ;
        RECT 162.240 35.600 162.410 35.810 ;
        RECT 163.620 35.600 163.790 35.810 ;
        RECT 165.455 35.650 165.575 35.760 ;
        RECT 165.920 35.600 166.090 35.790 ;
        RECT 170.520 35.620 170.690 35.810 ;
        RECT 171.255 35.620 171.425 35.810 ;
        RECT 175.855 35.620 176.025 35.810 ;
        RECT 178.340 35.600 178.510 35.790 ;
        RECT 179.730 35.655 179.890 35.765 ;
        RECT 180.640 35.620 180.810 35.810 ;
        RECT 184.320 35.620 184.490 35.810 ;
        RECT 187.540 35.600 187.710 35.790 ;
        RECT 188.460 35.600 188.630 35.790 ;
        RECT 196.740 35.620 196.910 35.810 ;
        RECT 197.200 35.620 197.370 35.810 ;
        RECT 200.880 35.600 201.050 35.790 ;
        RECT 201.340 35.600 201.510 35.810 ;
        RECT 204.095 35.650 204.215 35.760 ;
        RECT 204.835 35.620 205.005 35.810 ;
        RECT 208.700 35.620 208.870 35.810 ;
        RECT 210.535 35.650 210.655 35.760 ;
        RECT 212.840 35.600 213.010 35.790 ;
        RECT 213.295 35.650 213.415 35.760 ;
        RECT 214.230 35.645 214.390 35.755 ;
        RECT 214.405 35.620 214.575 35.810 ;
        RECT 215.415 35.620 215.585 35.810 ;
        RECT 222.500 35.620 222.670 35.810 ;
        RECT 223.880 35.600 224.050 35.790 ;
        RECT 224.340 35.600 224.510 35.790 ;
        RECT 226.180 35.620 226.350 35.810 ;
        RECT 227.100 35.620 227.270 35.810 ;
        RECT 228.940 35.620 229.110 35.810 ;
        RECT 233.540 35.600 233.710 35.790 ;
        RECT 237.220 35.600 237.390 35.790 ;
        RECT 237.680 35.600 237.850 35.790 ;
        RECT 238.600 35.620 238.770 35.810 ;
        RECT 239.980 35.760 240.150 35.810 ;
        RECT 239.975 35.650 240.150 35.760 ;
        RECT 239.980 35.620 240.150 35.650 ;
        RECT 240.440 35.600 240.610 35.790 ;
        RECT 249.180 35.620 249.350 35.810 ;
        RECT 249.640 35.600 249.810 35.790 ;
        RECT 251.935 35.650 252.055 35.760 ;
        RECT 252.860 35.620 253.030 35.810 ;
        RECT 253.330 35.645 253.490 35.755 ;
        RECT 254.240 35.600 254.410 35.810 ;
        RECT 265.280 35.790 265.445 35.810 ;
        RECT 267.580 35.790 267.730 35.810 ;
        RECT 263.440 35.600 263.610 35.790 ;
        RECT 265.280 35.620 265.450 35.790 ;
        RECT 265.740 35.600 265.910 35.790 ;
        RECT 267.580 35.620 267.750 35.790 ;
        RECT 268.050 35.655 268.210 35.765 ;
        RECT 268.960 35.620 269.130 35.810 ;
        RECT 271.255 35.650 271.375 35.760 ;
        RECT 271.720 35.600 271.890 35.790 ;
        RECT 278.625 35.620 278.795 35.840 ;
        RECT 280.755 35.810 281.690 35.840 ;
        RECT 281.700 35.810 287.210 36.620 ;
        RECT 287.220 35.810 292.730 36.620 ;
        RECT 292.740 35.810 298.250 36.620 ;
        RECT 298.260 35.810 303.770 36.620 ;
        RECT 303.790 35.895 304.220 36.680 ;
        RECT 304.240 35.810 307.910 36.620 ;
        RECT 307.920 35.810 309.750 36.490 ;
        RECT 309.760 35.810 311.130 36.620 ;
        RECT 280.920 35.600 281.090 35.790 ;
        RECT 281.840 35.620 282.010 35.810 ;
        RECT 286.440 35.600 286.610 35.790 ;
        RECT 287.360 35.620 287.530 35.810 ;
        RECT 290.130 35.645 290.290 35.755 ;
        RECT 291.500 35.600 291.670 35.790 ;
        RECT 292.880 35.620 293.050 35.810 ;
        RECT 297.020 35.600 297.190 35.790 ;
        RECT 298.400 35.620 298.570 35.810 ;
        RECT 302.540 35.600 302.710 35.790 ;
        RECT 304.380 35.620 304.550 35.810 ;
        RECT 308.060 35.600 308.230 35.790 ;
        RECT 309.440 35.620 309.610 35.810 ;
        RECT 310.820 35.600 310.990 35.810 ;
        RECT 162.100 34.790 163.470 35.600 ;
        RECT 163.480 34.790 165.310 35.600 ;
        RECT 165.780 34.920 174.970 35.600 ;
        RECT 170.290 34.700 171.220 34.920 ;
        RECT 174.050 34.690 174.970 34.920 ;
        RECT 175.075 34.920 178.540 35.600 ;
        RECT 178.660 34.920 187.850 35.600 ;
        RECT 175.075 34.690 175.995 34.920 ;
        RECT 178.660 34.690 179.580 34.920 ;
        RECT 182.410 34.700 183.340 34.920 ;
        RECT 187.870 34.730 188.300 35.515 ;
        RECT 188.320 34.920 197.510 35.600 ;
        RECT 192.830 34.700 193.760 34.920 ;
        RECT 196.590 34.690 197.510 34.920 ;
        RECT 197.615 34.920 201.080 35.600 ;
        RECT 201.200 34.920 210.390 35.600 ;
        RECT 210.410 34.920 213.150 35.600 ;
        RECT 197.615 34.690 198.535 34.920 ;
        RECT 205.710 34.700 206.640 34.920 ;
        RECT 209.470 34.690 210.390 34.920 ;
        RECT 213.630 34.730 214.060 35.515 ;
        RECT 215.000 34.920 224.190 35.600 ;
        RECT 224.200 34.920 233.390 35.600 ;
        RECT 215.000 34.690 215.920 34.920 ;
        RECT 218.750 34.700 219.680 34.920 ;
        RECT 228.710 34.700 229.640 34.920 ;
        RECT 232.470 34.690 233.390 34.920 ;
        RECT 233.400 34.790 234.770 35.600 ;
        RECT 234.790 34.920 237.530 35.600 ;
        RECT 237.540 34.790 239.370 35.600 ;
        RECT 239.390 34.730 239.820 35.515 ;
        RECT 240.300 34.920 249.490 35.600 ;
        RECT 244.810 34.700 245.740 34.920 ;
        RECT 248.570 34.690 249.490 34.920 ;
        RECT 249.500 34.790 253.170 35.600 ;
        RECT 254.100 34.920 263.290 35.600 ;
        RECT 258.610 34.700 259.540 34.920 ;
        RECT 262.370 34.690 263.290 34.920 ;
        RECT 263.300 34.790 265.130 35.600 ;
        RECT 265.150 34.730 265.580 35.515 ;
        RECT 265.600 34.790 271.110 35.600 ;
        RECT 271.580 34.920 280.770 35.600 ;
        RECT 276.090 34.700 277.020 34.920 ;
        RECT 279.850 34.690 280.770 34.920 ;
        RECT 280.780 34.790 286.290 35.600 ;
        RECT 286.300 34.790 289.970 35.600 ;
        RECT 290.910 34.730 291.340 35.515 ;
        RECT 291.360 34.790 296.870 35.600 ;
        RECT 296.880 34.790 302.390 35.600 ;
        RECT 302.400 34.790 307.910 35.600 ;
        RECT 307.920 34.790 309.750 35.600 ;
        RECT 309.760 34.790 311.130 35.600 ;
      LAYER nwell ;
        RECT 161.905 31.570 311.325 34.400 ;
      LAYER pwell ;
        RECT 162.100 30.370 163.470 31.180 ;
        RECT 163.480 30.370 165.310 31.180 ;
        RECT 170.290 31.050 171.220 31.270 ;
        RECT 174.050 31.050 174.970 31.280 ;
        RECT 165.780 30.370 174.970 31.050 ;
        RECT 174.990 30.455 175.420 31.240 ;
        RECT 175.440 31.050 176.370 31.280 ;
        RECT 175.440 30.370 179.340 31.050 ;
        RECT 179.580 30.370 182.330 31.180 ;
        RECT 182.340 31.050 183.260 31.280 ;
        RECT 186.090 31.050 187.020 31.270 ;
        RECT 194.740 31.050 195.670 31.280 ;
        RECT 182.340 30.370 191.530 31.050 ;
        RECT 191.770 30.370 195.670 31.050 ;
        RECT 195.680 30.370 197.050 31.180 ;
        RECT 199.715 31.050 200.635 31.280 ;
        RECT 197.170 30.370 200.635 31.050 ;
        RECT 200.750 30.455 201.180 31.240 ;
        RECT 201.200 31.050 202.130 31.280 ;
        RECT 201.200 30.370 205.100 31.050 ;
        RECT 205.340 30.370 207.170 31.180 ;
        RECT 207.180 31.050 208.100 31.280 ;
        RECT 210.930 31.050 211.860 31.270 ;
        RECT 216.475 31.050 217.395 31.280 ;
        RECT 207.180 30.370 216.370 31.050 ;
        RECT 216.475 30.370 219.940 31.050 ;
        RECT 220.060 30.370 225.570 31.180 ;
        RECT 226.510 30.455 226.940 31.240 ;
        RECT 226.960 31.050 227.890 31.280 ;
        RECT 234.675 31.050 235.595 31.280 ;
        RECT 226.960 30.370 230.860 31.050 ;
        RECT 232.130 30.370 235.595 31.050 ;
        RECT 235.700 31.050 236.620 31.280 ;
        RECT 239.450 31.050 240.380 31.270 ;
        RECT 235.700 30.370 244.890 31.050 ;
        RECT 244.900 30.370 250.410 31.180 ;
        RECT 250.420 30.370 252.250 31.180 ;
        RECT 252.270 30.455 252.700 31.240 ;
        RECT 252.720 30.370 258.230 31.180 ;
        RECT 258.720 30.370 260.070 31.280 ;
        RECT 260.080 30.370 265.590 31.180 ;
        RECT 265.600 30.370 271.110 31.180 ;
        RECT 271.120 30.370 276.630 31.180 ;
        RECT 276.640 30.370 278.010 31.180 ;
        RECT 278.030 30.455 278.460 31.240 ;
        RECT 278.480 30.370 283.990 31.180 ;
        RECT 284.000 30.370 289.510 31.180 ;
        RECT 289.520 30.370 295.030 31.180 ;
        RECT 295.040 30.370 300.550 31.180 ;
        RECT 300.560 30.370 303.310 31.180 ;
        RECT 303.790 30.455 304.220 31.240 ;
        RECT 304.240 30.370 309.750 31.180 ;
        RECT 309.760 30.370 311.130 31.180 ;
        RECT 162.240 30.160 162.410 30.370 ;
        RECT 163.620 30.180 163.790 30.370 ;
        RECT 165.000 30.160 165.170 30.350 ;
        RECT 165.460 30.320 165.630 30.350 ;
        RECT 165.455 30.210 165.630 30.320 ;
        RECT 165.460 30.160 165.630 30.210 ;
        RECT 165.920 30.180 166.090 30.370 ;
        RECT 168.215 30.210 168.335 30.320 ;
        RECT 171.900 30.160 172.070 30.350 ;
        RECT 172.635 30.160 172.805 30.350 ;
        RECT 175.855 30.180 176.025 30.370 ;
        RECT 176.500 30.160 176.670 30.350 ;
        RECT 179.720 30.180 179.890 30.370 ;
        RECT 180.180 30.160 180.350 30.350 ;
        RECT 184.135 30.160 184.305 30.350 ;
        RECT 188.735 30.160 188.905 30.350 ;
        RECT 191.220 30.180 191.390 30.370 ;
        RECT 192.595 30.210 192.715 30.320 ;
        RECT 195.085 30.180 195.255 30.370 ;
        RECT 195.820 30.180 195.990 30.370 ;
        RECT 196.280 30.160 196.450 30.350 ;
        RECT 197.200 30.180 197.370 30.370 ;
        RECT 201.615 30.180 201.785 30.370 ;
        RECT 205.480 30.160 205.650 30.370 ;
        RECT 205.940 30.160 206.110 30.350 ;
        RECT 211.920 30.160 212.090 30.350 ;
        RECT 212.380 30.160 212.550 30.350 ;
        RECT 214.220 30.160 214.390 30.350 ;
        RECT 216.060 30.180 216.230 30.370 ;
        RECT 219.740 30.160 219.910 30.370 ;
        RECT 220.200 30.180 220.370 30.370 ;
        RECT 225.260 30.160 225.430 30.350 ;
        RECT 225.730 30.215 225.890 30.325 ;
        RECT 227.375 30.180 227.545 30.370 ;
        RECT 230.780 30.160 230.950 30.350 ;
        RECT 231.250 30.215 231.410 30.325 ;
        RECT 232.160 30.180 232.330 30.370 ;
        RECT 236.300 30.160 236.470 30.350 ;
        RECT 239.055 30.210 239.175 30.320 ;
        RECT 239.980 30.160 240.150 30.350 ;
        RECT 244.580 30.180 244.750 30.370 ;
        RECT 245.040 30.180 245.210 30.370 ;
        RECT 245.500 30.160 245.670 30.350 ;
        RECT 250.560 30.180 250.730 30.370 ;
        RECT 251.020 30.160 251.190 30.350 ;
        RECT 252.860 30.180 253.030 30.370 ;
        RECT 256.540 30.160 256.710 30.350 ;
        RECT 258.375 30.210 258.495 30.320 ;
        RECT 259.755 30.180 259.925 30.370 ;
        RECT 260.220 30.180 260.390 30.370 ;
        RECT 262.060 30.160 262.230 30.350 ;
        RECT 264.815 30.210 264.935 30.320 ;
        RECT 265.740 30.160 265.910 30.370 ;
        RECT 271.260 30.160 271.430 30.370 ;
        RECT 276.780 30.160 276.950 30.370 ;
        RECT 278.620 30.180 278.790 30.370 ;
        RECT 282.300 30.160 282.470 30.350 ;
        RECT 284.140 30.180 284.310 30.370 ;
        RECT 287.820 30.160 287.990 30.350 ;
        RECT 289.660 30.180 289.830 30.370 ;
        RECT 290.575 30.210 290.695 30.320 ;
        RECT 291.500 30.160 291.670 30.350 ;
        RECT 295.180 30.180 295.350 30.370 ;
        RECT 297.020 30.160 297.190 30.350 ;
        RECT 300.700 30.180 300.870 30.370 ;
        RECT 302.540 30.160 302.710 30.350 ;
        RECT 303.455 30.210 303.575 30.320 ;
        RECT 304.380 30.180 304.550 30.370 ;
        RECT 308.060 30.160 308.230 30.350 ;
        RECT 310.820 30.160 310.990 30.370 ;
        RECT 162.100 29.350 163.470 30.160 ;
        RECT 163.480 29.480 165.310 30.160 ;
        RECT 163.480 29.250 164.825 29.480 ;
        RECT 165.320 29.350 168.070 30.160 ;
        RECT 168.635 29.480 172.100 30.160 ;
        RECT 172.220 29.480 176.120 30.160 ;
        RECT 176.470 29.480 179.935 30.160 ;
        RECT 180.150 29.480 183.615 30.160 ;
        RECT 168.635 29.250 169.555 29.480 ;
        RECT 172.220 29.250 173.150 29.480 ;
        RECT 179.015 29.250 179.935 29.480 ;
        RECT 182.695 29.250 183.615 29.480 ;
        RECT 183.720 29.480 187.620 30.160 ;
        RECT 183.720 29.250 184.650 29.480 ;
        RECT 187.870 29.290 188.300 30.075 ;
        RECT 188.320 29.480 192.220 30.160 ;
        RECT 193.015 29.480 196.480 30.160 ;
        RECT 196.600 29.480 205.790 30.160 ;
        RECT 188.320 29.250 189.250 29.480 ;
        RECT 193.015 29.250 193.935 29.480 ;
        RECT 196.600 29.250 197.520 29.480 ;
        RECT 200.350 29.260 201.280 29.480 ;
        RECT 205.800 29.350 208.550 30.160 ;
        RECT 208.655 29.480 212.120 30.160 ;
        RECT 208.655 29.250 209.575 29.480 ;
        RECT 212.240 29.350 213.610 30.160 ;
        RECT 213.630 29.290 214.060 30.075 ;
        RECT 214.080 29.350 219.590 30.160 ;
        RECT 219.600 29.350 225.110 30.160 ;
        RECT 225.120 29.350 230.630 30.160 ;
        RECT 230.640 29.350 236.150 30.160 ;
        RECT 236.160 29.350 238.910 30.160 ;
        RECT 239.390 29.290 239.820 30.075 ;
        RECT 239.840 29.350 245.350 30.160 ;
        RECT 245.360 29.350 250.870 30.160 ;
        RECT 250.880 29.350 256.390 30.160 ;
        RECT 256.400 29.350 261.910 30.160 ;
        RECT 261.920 29.350 264.670 30.160 ;
        RECT 265.150 29.290 265.580 30.075 ;
        RECT 265.600 29.350 271.110 30.160 ;
        RECT 271.120 29.350 276.630 30.160 ;
        RECT 276.640 29.350 282.150 30.160 ;
        RECT 282.160 29.350 287.670 30.160 ;
        RECT 287.680 29.350 290.430 30.160 ;
        RECT 290.910 29.290 291.340 30.075 ;
        RECT 291.360 29.350 296.870 30.160 ;
        RECT 296.880 29.350 302.390 30.160 ;
        RECT 302.400 29.350 307.910 30.160 ;
        RECT 307.920 29.350 309.750 30.160 ;
        RECT 309.760 29.350 311.130 30.160 ;
      LAYER nwell ;
        RECT 161.905 26.130 311.325 28.960 ;
      LAYER pwell ;
        RECT 162.100 24.930 163.470 25.740 ;
        RECT 163.480 24.930 168.990 25.740 ;
        RECT 169.000 24.930 170.830 25.740 ;
        RECT 171.395 25.610 172.315 25.840 ;
        RECT 171.395 24.930 174.860 25.610 ;
        RECT 174.990 25.015 175.420 25.800 ;
        RECT 175.535 25.610 176.455 25.840 ;
        RECT 175.535 24.930 179.000 25.610 ;
        RECT 179.120 24.930 184.630 25.740 ;
        RECT 184.640 24.930 188.310 25.740 ;
        RECT 191.895 25.610 192.815 25.840 ;
        RECT 189.350 24.930 192.815 25.610 ;
        RECT 192.920 24.930 196.590 25.740 ;
        RECT 196.600 24.930 197.970 25.740 ;
        RECT 197.990 24.930 200.730 25.610 ;
        RECT 200.750 25.015 201.180 25.800 ;
        RECT 201.200 24.930 204.870 25.740 ;
        RECT 207.995 25.610 208.915 25.840 ;
        RECT 205.450 24.930 208.915 25.610 ;
        RECT 209.020 24.930 214.530 25.740 ;
        RECT 214.540 24.930 220.050 25.740 ;
        RECT 220.060 24.930 225.570 25.740 ;
        RECT 226.510 25.015 226.940 25.800 ;
        RECT 226.960 24.930 232.470 25.740 ;
        RECT 232.480 24.930 237.990 25.740 ;
        RECT 238.000 24.930 243.510 25.740 ;
        RECT 243.520 24.930 249.030 25.740 ;
        RECT 249.040 24.930 251.790 25.740 ;
        RECT 252.270 25.015 252.700 25.800 ;
        RECT 252.720 24.930 258.230 25.740 ;
        RECT 258.240 24.930 263.750 25.740 ;
        RECT 263.760 24.930 269.270 25.740 ;
        RECT 269.280 24.930 274.790 25.740 ;
        RECT 274.800 24.930 277.550 25.740 ;
        RECT 278.030 25.015 278.460 25.800 ;
        RECT 278.480 24.930 283.990 25.740 ;
        RECT 284.000 24.930 289.510 25.740 ;
        RECT 289.520 24.930 295.030 25.740 ;
        RECT 295.040 24.930 300.550 25.740 ;
        RECT 300.560 24.930 303.310 25.740 ;
        RECT 303.790 25.015 304.220 25.800 ;
        RECT 304.240 24.930 309.750 25.740 ;
        RECT 309.760 24.930 311.130 25.740 ;
        RECT 162.240 24.720 162.410 24.930 ;
        RECT 163.620 24.720 163.790 24.930 ;
        RECT 169.140 24.720 169.310 24.930 ;
        RECT 170.975 24.770 171.095 24.880 ;
        RECT 174.660 24.720 174.830 24.930 ;
        RECT 178.800 24.740 178.970 24.930 ;
        RECT 179.260 24.740 179.430 24.930 ;
        RECT 180.180 24.720 180.350 24.910 ;
        RECT 184.780 24.740 184.950 24.930 ;
        RECT 185.700 24.720 185.870 24.910 ;
        RECT 187.535 24.770 187.655 24.880 ;
        RECT 188.460 24.720 188.630 24.910 ;
        RECT 189.380 24.740 189.550 24.930 ;
        RECT 193.060 24.740 193.230 24.930 ;
        RECT 193.980 24.720 194.150 24.910 ;
        RECT 196.740 24.740 196.910 24.930 ;
        RECT 199.500 24.720 199.670 24.910 ;
        RECT 200.420 24.740 200.590 24.930 ;
        RECT 201.340 24.740 201.510 24.930 ;
        RECT 205.020 24.880 205.190 24.910 ;
        RECT 205.015 24.770 205.190 24.880 ;
        RECT 205.020 24.720 205.190 24.770 ;
        RECT 205.480 24.740 205.650 24.930 ;
        RECT 209.160 24.740 209.330 24.930 ;
        RECT 210.540 24.720 210.710 24.910 ;
        RECT 213.295 24.770 213.415 24.880 ;
        RECT 214.220 24.720 214.390 24.910 ;
        RECT 214.680 24.740 214.850 24.930 ;
        RECT 219.740 24.720 219.910 24.910 ;
        RECT 220.200 24.740 220.370 24.930 ;
        RECT 225.260 24.720 225.430 24.910 ;
        RECT 225.730 24.775 225.890 24.885 ;
        RECT 227.100 24.740 227.270 24.930 ;
        RECT 230.780 24.720 230.950 24.910 ;
        RECT 232.620 24.740 232.790 24.930 ;
        RECT 236.300 24.720 236.470 24.910 ;
        RECT 238.140 24.740 238.310 24.930 ;
        RECT 239.055 24.770 239.175 24.880 ;
        RECT 239.980 24.720 240.150 24.910 ;
        RECT 243.660 24.740 243.830 24.930 ;
        RECT 245.500 24.720 245.670 24.910 ;
        RECT 249.180 24.740 249.350 24.930 ;
        RECT 251.020 24.720 251.190 24.910 ;
        RECT 251.935 24.770 252.055 24.880 ;
        RECT 252.860 24.740 253.030 24.930 ;
        RECT 256.540 24.720 256.710 24.910 ;
        RECT 258.380 24.740 258.550 24.930 ;
        RECT 262.060 24.720 262.230 24.910 ;
        RECT 263.900 24.740 264.070 24.930 ;
        RECT 264.815 24.770 264.935 24.880 ;
        RECT 265.740 24.720 265.910 24.910 ;
        RECT 269.420 24.740 269.590 24.930 ;
        RECT 271.260 24.720 271.430 24.910 ;
        RECT 274.940 24.740 275.110 24.930 ;
        RECT 276.780 24.720 276.950 24.910 ;
        RECT 277.695 24.770 277.815 24.880 ;
        RECT 278.620 24.740 278.790 24.930 ;
        RECT 282.300 24.720 282.470 24.910 ;
        RECT 284.140 24.740 284.310 24.930 ;
        RECT 287.820 24.720 287.990 24.910 ;
        RECT 289.660 24.740 289.830 24.930 ;
        RECT 290.575 24.770 290.695 24.880 ;
        RECT 291.500 24.720 291.670 24.910 ;
        RECT 295.180 24.740 295.350 24.930 ;
        RECT 297.020 24.720 297.190 24.910 ;
        RECT 300.700 24.740 300.870 24.930 ;
        RECT 302.540 24.720 302.710 24.910 ;
        RECT 303.455 24.770 303.575 24.880 ;
        RECT 304.380 24.740 304.550 24.930 ;
        RECT 308.060 24.720 308.230 24.910 ;
        RECT 310.820 24.720 310.990 24.930 ;
        RECT 162.100 23.910 163.470 24.720 ;
        RECT 163.480 23.910 168.990 24.720 ;
        RECT 169.000 23.910 174.510 24.720 ;
        RECT 174.520 23.910 180.030 24.720 ;
        RECT 180.040 23.910 185.550 24.720 ;
        RECT 185.560 23.910 187.390 24.720 ;
        RECT 187.870 23.850 188.300 24.635 ;
        RECT 188.320 23.910 193.830 24.720 ;
        RECT 193.840 23.910 199.350 24.720 ;
        RECT 199.360 23.910 204.870 24.720 ;
        RECT 204.880 23.910 210.390 24.720 ;
        RECT 210.400 23.910 213.150 24.720 ;
        RECT 213.630 23.850 214.060 24.635 ;
        RECT 214.080 23.910 219.590 24.720 ;
        RECT 219.600 23.910 225.110 24.720 ;
        RECT 225.120 23.910 230.630 24.720 ;
        RECT 230.640 23.910 236.150 24.720 ;
        RECT 236.160 23.910 238.910 24.720 ;
        RECT 239.390 23.850 239.820 24.635 ;
        RECT 239.840 23.910 245.350 24.720 ;
        RECT 245.360 23.910 250.870 24.720 ;
        RECT 250.880 23.910 256.390 24.720 ;
        RECT 256.400 23.910 261.910 24.720 ;
        RECT 261.920 23.910 264.670 24.720 ;
        RECT 265.150 23.850 265.580 24.635 ;
        RECT 265.600 23.910 271.110 24.720 ;
        RECT 271.120 23.910 276.630 24.720 ;
        RECT 276.640 23.910 282.150 24.720 ;
        RECT 282.160 23.910 287.670 24.720 ;
        RECT 287.680 23.910 290.430 24.720 ;
        RECT 290.910 23.850 291.340 24.635 ;
        RECT 291.360 23.910 296.870 24.720 ;
        RECT 296.880 23.910 302.390 24.720 ;
        RECT 302.400 23.910 307.910 24.720 ;
        RECT 307.920 23.910 309.750 24.720 ;
        RECT 309.760 23.910 311.130 24.720 ;
      LAYER nwell ;
        RECT 161.905 20.690 311.325 23.520 ;
      LAYER pwell ;
        RECT 162.100 19.490 163.470 20.300 ;
        RECT 163.480 19.490 168.990 20.300 ;
        RECT 169.000 19.490 174.510 20.300 ;
        RECT 174.990 19.575 175.420 20.360 ;
        RECT 175.440 19.490 180.950 20.300 ;
        RECT 180.960 19.490 186.470 20.300 ;
        RECT 186.480 19.490 191.990 20.300 ;
        RECT 192.000 19.490 197.510 20.300 ;
        RECT 197.520 19.490 200.270 20.300 ;
        RECT 200.750 19.575 201.180 20.360 ;
        RECT 201.200 19.490 206.710 20.300 ;
        RECT 206.720 19.490 212.230 20.300 ;
        RECT 212.240 19.490 217.750 20.300 ;
        RECT 217.760 19.490 223.270 20.300 ;
        RECT 223.280 19.490 226.030 20.300 ;
        RECT 226.510 19.575 226.940 20.360 ;
        RECT 226.960 19.490 232.470 20.300 ;
        RECT 232.480 19.490 237.990 20.300 ;
        RECT 238.000 19.490 243.510 20.300 ;
        RECT 243.520 19.490 249.030 20.300 ;
        RECT 249.040 19.490 251.790 20.300 ;
        RECT 252.270 19.575 252.700 20.360 ;
        RECT 252.720 19.490 258.230 20.300 ;
        RECT 258.240 19.490 263.750 20.300 ;
        RECT 263.760 19.490 269.270 20.300 ;
        RECT 269.280 19.490 274.790 20.300 ;
        RECT 274.800 19.490 277.550 20.300 ;
        RECT 278.030 19.575 278.460 20.360 ;
        RECT 278.480 19.490 283.990 20.300 ;
        RECT 284.000 19.490 289.510 20.300 ;
        RECT 289.520 19.490 295.030 20.300 ;
        RECT 295.040 19.490 300.550 20.300 ;
        RECT 300.560 19.490 303.310 20.300 ;
        RECT 303.790 19.575 304.220 20.360 ;
        RECT 304.240 19.490 309.750 20.300 ;
        RECT 309.760 19.490 311.130 20.300 ;
        RECT 162.240 19.280 162.410 19.490 ;
        RECT 163.620 19.280 163.790 19.490 ;
        RECT 169.140 19.280 169.310 19.490 ;
        RECT 174.660 19.440 174.830 19.470 ;
        RECT 174.655 19.330 174.830 19.440 ;
        RECT 174.660 19.280 174.830 19.330 ;
        RECT 175.580 19.300 175.750 19.490 ;
        RECT 180.180 19.280 180.350 19.470 ;
        RECT 181.100 19.300 181.270 19.490 ;
        RECT 185.700 19.280 185.870 19.470 ;
        RECT 186.620 19.300 186.790 19.490 ;
        RECT 187.535 19.330 187.655 19.440 ;
        RECT 188.460 19.280 188.630 19.470 ;
        RECT 192.140 19.300 192.310 19.490 ;
        RECT 193.980 19.280 194.150 19.470 ;
        RECT 197.660 19.300 197.830 19.490 ;
        RECT 199.500 19.280 199.670 19.470 ;
        RECT 200.415 19.330 200.535 19.440 ;
        RECT 201.340 19.300 201.510 19.490 ;
        RECT 205.020 19.280 205.190 19.470 ;
        RECT 206.860 19.300 207.030 19.490 ;
        RECT 210.540 19.280 210.710 19.470 ;
        RECT 212.380 19.300 212.550 19.490 ;
        RECT 213.295 19.330 213.415 19.440 ;
        RECT 214.220 19.280 214.390 19.470 ;
        RECT 217.900 19.300 218.070 19.490 ;
        RECT 219.740 19.280 219.910 19.470 ;
        RECT 223.420 19.300 223.590 19.490 ;
        RECT 225.260 19.280 225.430 19.470 ;
        RECT 226.175 19.330 226.295 19.440 ;
        RECT 227.100 19.300 227.270 19.490 ;
        RECT 230.780 19.280 230.950 19.470 ;
        RECT 232.620 19.300 232.790 19.490 ;
        RECT 236.300 19.280 236.470 19.470 ;
        RECT 238.140 19.300 238.310 19.490 ;
        RECT 239.055 19.330 239.175 19.440 ;
        RECT 239.980 19.280 240.150 19.470 ;
        RECT 243.660 19.300 243.830 19.490 ;
        RECT 245.500 19.280 245.670 19.470 ;
        RECT 249.180 19.300 249.350 19.490 ;
        RECT 251.020 19.280 251.190 19.470 ;
        RECT 251.935 19.330 252.055 19.440 ;
        RECT 252.860 19.300 253.030 19.490 ;
        RECT 256.540 19.280 256.710 19.470 ;
        RECT 258.380 19.300 258.550 19.490 ;
        RECT 262.060 19.280 262.230 19.470 ;
        RECT 263.900 19.300 264.070 19.490 ;
        RECT 264.815 19.330 264.935 19.440 ;
        RECT 265.740 19.280 265.910 19.470 ;
        RECT 269.420 19.300 269.590 19.490 ;
        RECT 271.260 19.280 271.430 19.470 ;
        RECT 274.940 19.300 275.110 19.490 ;
        RECT 276.780 19.280 276.950 19.470 ;
        RECT 277.695 19.330 277.815 19.440 ;
        RECT 278.620 19.300 278.790 19.490 ;
        RECT 282.300 19.280 282.470 19.470 ;
        RECT 284.140 19.300 284.310 19.490 ;
        RECT 287.820 19.280 287.990 19.470 ;
        RECT 289.660 19.300 289.830 19.490 ;
        RECT 290.575 19.330 290.695 19.440 ;
        RECT 291.500 19.280 291.670 19.470 ;
        RECT 295.180 19.300 295.350 19.490 ;
        RECT 297.020 19.280 297.190 19.470 ;
        RECT 300.700 19.300 300.870 19.490 ;
        RECT 302.540 19.280 302.710 19.470 ;
        RECT 303.455 19.330 303.575 19.440 ;
        RECT 304.380 19.300 304.550 19.490 ;
        RECT 308.060 19.280 308.230 19.470 ;
        RECT 310.820 19.280 310.990 19.490 ;
        RECT 162.100 18.470 163.470 19.280 ;
        RECT 163.480 18.470 168.990 19.280 ;
        RECT 169.000 18.470 174.510 19.280 ;
        RECT 174.520 18.470 180.030 19.280 ;
        RECT 180.040 18.470 185.550 19.280 ;
        RECT 185.560 18.470 187.390 19.280 ;
        RECT 187.870 18.410 188.300 19.195 ;
        RECT 188.320 18.470 193.830 19.280 ;
        RECT 193.840 18.470 199.350 19.280 ;
        RECT 199.360 18.470 204.870 19.280 ;
        RECT 204.880 18.470 210.390 19.280 ;
        RECT 210.400 18.470 213.150 19.280 ;
        RECT 213.630 18.410 214.060 19.195 ;
        RECT 214.080 18.470 219.590 19.280 ;
        RECT 219.600 18.470 225.110 19.280 ;
        RECT 225.120 18.470 230.630 19.280 ;
        RECT 230.640 18.470 236.150 19.280 ;
        RECT 236.160 18.470 238.910 19.280 ;
        RECT 239.390 18.410 239.820 19.195 ;
        RECT 239.840 18.470 245.350 19.280 ;
        RECT 245.360 18.470 250.870 19.280 ;
        RECT 250.880 18.470 256.390 19.280 ;
        RECT 256.400 18.470 261.910 19.280 ;
        RECT 261.920 18.470 264.670 19.280 ;
        RECT 265.150 18.410 265.580 19.195 ;
        RECT 265.600 18.470 271.110 19.280 ;
        RECT 271.120 18.470 276.630 19.280 ;
        RECT 276.640 18.470 282.150 19.280 ;
        RECT 282.160 18.470 287.670 19.280 ;
        RECT 287.680 18.470 290.430 19.280 ;
        RECT 290.910 18.410 291.340 19.195 ;
        RECT 291.360 18.470 296.870 19.280 ;
        RECT 296.880 18.470 302.390 19.280 ;
        RECT 302.400 18.470 307.910 19.280 ;
        RECT 307.920 18.470 309.750 19.280 ;
        RECT 309.760 18.470 311.130 19.280 ;
      LAYER nwell ;
        RECT 161.905 15.250 311.325 18.080 ;
      LAYER pwell ;
        RECT 162.100 14.050 163.470 14.860 ;
        RECT 163.480 14.050 168.990 14.860 ;
        RECT 169.000 14.050 174.510 14.860 ;
        RECT 174.990 14.135 175.420 14.920 ;
        RECT 175.440 14.050 180.950 14.860 ;
        RECT 180.960 14.050 186.470 14.860 ;
        RECT 186.480 14.050 187.850 14.860 ;
        RECT 187.870 14.135 188.300 14.920 ;
        RECT 188.320 14.050 193.830 14.860 ;
        RECT 193.840 14.050 199.350 14.860 ;
        RECT 199.360 14.050 200.730 14.860 ;
        RECT 200.750 14.135 201.180 14.920 ;
        RECT 201.200 14.050 206.710 14.860 ;
        RECT 206.720 14.050 212.230 14.860 ;
        RECT 212.240 14.050 213.610 14.860 ;
        RECT 213.630 14.135 214.060 14.920 ;
        RECT 214.080 14.050 219.590 14.860 ;
        RECT 219.600 14.050 225.110 14.860 ;
        RECT 225.120 14.050 226.490 14.860 ;
        RECT 226.510 14.135 226.940 14.920 ;
        RECT 226.960 14.050 232.470 14.860 ;
        RECT 232.480 14.050 237.990 14.860 ;
        RECT 238.000 14.050 239.370 14.860 ;
        RECT 239.390 14.135 239.820 14.920 ;
        RECT 239.840 14.050 245.350 14.860 ;
        RECT 245.360 14.050 250.870 14.860 ;
        RECT 250.880 14.050 252.250 14.860 ;
        RECT 252.270 14.135 252.700 14.920 ;
        RECT 252.720 14.050 258.230 14.860 ;
        RECT 258.240 14.050 263.750 14.860 ;
        RECT 263.760 14.050 265.130 14.860 ;
        RECT 265.150 14.135 265.580 14.920 ;
        RECT 265.600 14.050 271.110 14.860 ;
        RECT 271.120 14.050 276.630 14.860 ;
        RECT 276.640 14.050 278.010 14.860 ;
        RECT 278.030 14.135 278.460 14.920 ;
        RECT 278.480 14.050 283.990 14.860 ;
        RECT 284.000 14.050 289.510 14.860 ;
        RECT 289.520 14.050 290.890 14.860 ;
        RECT 290.910 14.135 291.340 14.920 ;
        RECT 291.360 14.050 296.870 14.860 ;
        RECT 296.880 14.050 302.390 14.860 ;
        RECT 302.400 14.050 303.770 14.860 ;
        RECT 303.790 14.135 304.220 14.920 ;
        RECT 304.240 14.050 309.750 14.860 ;
        RECT 309.760 14.050 311.130 14.860 ;
        RECT 162.240 13.860 162.410 14.050 ;
        RECT 163.620 13.860 163.790 14.050 ;
        RECT 169.140 13.860 169.310 14.050 ;
        RECT 174.655 13.890 174.775 14.000 ;
        RECT 175.580 13.860 175.750 14.050 ;
        RECT 181.100 13.860 181.270 14.050 ;
        RECT 186.620 13.860 186.790 14.050 ;
        RECT 188.460 13.860 188.630 14.050 ;
        RECT 193.980 13.860 194.150 14.050 ;
        RECT 199.500 13.860 199.670 14.050 ;
        RECT 201.340 13.860 201.510 14.050 ;
        RECT 206.860 13.860 207.030 14.050 ;
        RECT 212.380 13.860 212.550 14.050 ;
        RECT 214.220 13.860 214.390 14.050 ;
        RECT 219.740 13.860 219.910 14.050 ;
        RECT 225.260 13.860 225.430 14.050 ;
        RECT 227.100 13.860 227.270 14.050 ;
        RECT 232.620 13.860 232.790 14.050 ;
        RECT 238.140 13.860 238.310 14.050 ;
        RECT 239.980 13.860 240.150 14.050 ;
        RECT 245.500 13.860 245.670 14.050 ;
        RECT 251.020 13.860 251.190 14.050 ;
        RECT 252.860 13.860 253.030 14.050 ;
        RECT 258.380 13.860 258.550 14.050 ;
        RECT 263.900 13.860 264.070 14.050 ;
        RECT 265.740 13.860 265.910 14.050 ;
        RECT 271.260 13.860 271.430 14.050 ;
        RECT 276.780 13.860 276.950 14.050 ;
        RECT 278.620 13.860 278.790 14.050 ;
        RECT 284.140 13.860 284.310 14.050 ;
        RECT 289.660 13.860 289.830 14.050 ;
        RECT 291.500 13.860 291.670 14.050 ;
        RECT 297.020 13.860 297.190 14.050 ;
        RECT 302.540 13.860 302.710 14.050 ;
        RECT 304.380 13.860 304.550 14.050 ;
        RECT 310.820 13.860 310.990 14.050 ;
      LAYER nwell ;
        RECT 3.250 3.250 156.750 5.750 ;
      LAYER li1 ;
        RECT 4.300 222.030 102.625 222.430 ;
        RECT 4.300 4.700 4.700 222.030 ;
        RECT 62.895 216.545 99.045 217.075 ;
        RECT 62.895 213.695 63.425 216.545 ;
        RECT 63.925 215.855 80.385 216.025 ;
        RECT 63.925 214.385 64.155 215.855 ;
        RECT 80.155 214.385 80.385 215.855 ;
        RECT 63.925 214.215 80.385 214.385 ;
        RECT 80.885 213.695 81.055 216.545 ;
        RECT 81.555 215.855 98.015 216.025 ;
        RECT 81.555 214.385 81.785 215.855 ;
        RECT 97.785 214.385 98.015 215.855 ;
        RECT 81.555 214.215 98.015 214.385 ;
        RECT 98.515 213.695 99.045 216.545 ;
        RECT 62.895 213.525 99.045 213.695 ;
        RECT 9.325 211.690 45.335 211.860 ;
        RECT 9.325 201.840 9.495 211.690 ;
        RECT 10.225 211.000 18.225 211.170 ;
        RECT 18.515 211.000 26.515 211.170 ;
        RECT 9.995 202.745 10.165 210.785 ;
        RECT 18.285 202.745 18.455 210.785 ;
        RECT 26.575 202.745 26.745 210.785 ;
        RECT 10.225 202.360 18.225 202.530 ;
        RECT 18.515 202.360 26.515 202.530 ;
        RECT 27.245 201.840 27.415 211.690 ;
        RECT 28.145 211.000 36.145 211.170 ;
        RECT 36.435 211.000 44.435 211.170 ;
        RECT 27.915 202.745 28.085 210.785 ;
        RECT 36.205 202.745 36.375 210.785 ;
        RECT 44.495 202.745 44.665 210.785 ;
        RECT 28.145 202.360 36.145 202.530 ;
        RECT 36.435 202.360 44.435 202.530 ;
        RECT 45.165 201.840 45.335 211.690 ;
        RECT 62.895 210.675 63.425 213.525 ;
        RECT 64.155 212.835 80.155 213.005 ;
        RECT 63.925 211.580 64.095 212.620 ;
        RECT 80.215 211.580 80.385 212.620 ;
        RECT 64.155 211.195 80.155 211.365 ;
        RECT 80.885 210.675 81.055 213.525 ;
        RECT 81.785 212.835 97.785 213.005 ;
        RECT 81.555 211.580 81.725 212.620 ;
        RECT 97.845 211.580 98.015 212.620 ;
        RECT 81.785 211.195 97.785 211.365 ;
        RECT 98.515 210.675 99.045 213.525 ;
        RECT 62.895 210.505 99.045 210.675 ;
        RECT 9.325 201.670 45.335 201.840 ;
        RECT 9.325 191.820 9.495 201.670 ;
        RECT 10.225 200.980 18.225 201.150 ;
        RECT 18.515 200.980 26.515 201.150 ;
        RECT 9.995 192.725 10.165 200.765 ;
        RECT 18.285 192.725 18.455 200.765 ;
        RECT 26.575 192.725 26.745 200.765 ;
        RECT 10.225 192.340 18.225 192.510 ;
        RECT 18.515 192.340 26.515 192.510 ;
        RECT 27.245 191.820 27.415 201.670 ;
        RECT 28.145 200.980 36.145 201.150 ;
        RECT 36.435 200.980 44.435 201.150 ;
        RECT 27.915 192.725 28.085 200.765 ;
        RECT 36.205 192.725 36.375 200.765 ;
        RECT 44.495 192.725 44.665 200.765 ;
        RECT 28.145 192.340 36.145 192.510 ;
        RECT 36.435 192.340 44.435 192.510 ;
        RECT 45.165 191.820 45.335 201.670 ;
        RECT 9.325 191.650 45.335 191.820 ;
        RECT 49.250 210.180 56.310 210.350 ;
        RECT 9.325 190.700 15.415 190.870 ;
        RECT 9.325 180.850 9.495 190.700 ;
        RECT 10.225 190.010 12.225 190.180 ;
        RECT 12.515 190.010 14.515 190.180 ;
        RECT 9.995 181.755 10.165 189.795 ;
        RECT 12.285 181.755 12.455 189.795 ;
        RECT 14.575 181.755 14.745 189.795 ;
        RECT 10.225 181.370 12.225 181.540 ;
        RECT 12.515 181.370 14.515 181.540 ;
        RECT 15.245 180.850 15.415 190.700 ;
        RECT 9.325 180.680 15.415 180.850 ;
        RECT 16.345 190.700 45.335 190.870 ;
        RECT 16.345 180.850 16.515 190.700 ;
        RECT 17.245 190.010 19.245 190.180 ;
        RECT 19.535 190.010 21.535 190.180 ;
        RECT 21.825 190.010 23.825 190.180 ;
        RECT 24.115 190.010 26.115 190.180 ;
        RECT 26.405 190.010 28.405 190.180 ;
        RECT 28.695 190.010 30.695 190.180 ;
        RECT 30.985 190.010 32.985 190.180 ;
        RECT 33.275 190.010 35.275 190.180 ;
        RECT 35.565 190.010 37.565 190.180 ;
        RECT 37.855 190.010 39.855 190.180 ;
        RECT 40.145 190.010 42.145 190.180 ;
        RECT 42.435 190.010 44.435 190.180 ;
        RECT 17.015 181.755 17.185 189.795 ;
        RECT 19.305 181.755 19.475 189.795 ;
        RECT 21.595 181.755 21.765 189.795 ;
        RECT 23.885 181.755 24.055 189.795 ;
        RECT 26.175 181.755 26.345 189.795 ;
        RECT 28.465 181.755 28.635 189.795 ;
        RECT 30.755 181.755 30.925 189.795 ;
        RECT 33.045 181.755 33.215 189.795 ;
        RECT 35.335 181.755 35.505 189.795 ;
        RECT 37.625 181.755 37.795 189.795 ;
        RECT 39.915 181.755 40.085 189.795 ;
        RECT 42.205 181.755 42.375 189.795 ;
        RECT 44.495 181.755 44.665 189.795 ;
        RECT 17.245 181.370 19.245 181.540 ;
        RECT 19.535 181.370 21.535 181.540 ;
        RECT 21.825 181.370 23.825 181.540 ;
        RECT 24.115 181.370 26.115 181.540 ;
        RECT 26.405 181.370 28.405 181.540 ;
        RECT 28.695 181.370 30.695 181.540 ;
        RECT 30.985 181.370 32.985 181.540 ;
        RECT 33.275 181.370 35.275 181.540 ;
        RECT 35.565 181.370 37.565 181.540 ;
        RECT 37.855 181.370 39.855 181.540 ;
        RECT 40.145 181.370 42.145 181.540 ;
        RECT 42.435 181.370 44.435 181.540 ;
        RECT 45.165 180.850 45.335 190.700 ;
        RECT 49.250 187.850 49.420 210.180 ;
        RECT 50.095 207.435 50.785 209.595 ;
        RECT 51.265 207.435 51.955 209.595 ;
        RECT 52.435 207.435 53.125 209.595 ;
        RECT 53.605 207.435 54.295 209.595 ;
        RECT 54.775 207.435 55.465 209.595 ;
        RECT 50.095 188.435 50.785 190.595 ;
        RECT 51.265 188.435 51.955 190.595 ;
        RECT 52.435 188.435 53.125 190.595 ;
        RECT 53.605 188.435 54.295 190.595 ;
        RECT 54.775 188.435 55.465 190.595 ;
        RECT 56.140 187.850 56.310 210.180 ;
        RECT 49.250 187.680 56.310 187.850 ;
        RECT 62.895 207.655 63.425 210.505 ;
        RECT 64.155 209.815 80.155 209.985 ;
        RECT 63.925 208.560 64.095 209.600 ;
        RECT 80.215 208.560 80.385 209.600 ;
        RECT 64.155 208.175 80.155 208.345 ;
        RECT 80.885 207.655 81.055 210.505 ;
        RECT 81.785 209.815 97.785 209.985 ;
        RECT 81.555 208.560 81.725 209.600 ;
        RECT 97.845 208.560 98.015 209.600 ;
        RECT 81.785 208.175 97.785 208.345 ;
        RECT 98.515 207.655 99.045 210.505 ;
        RECT 62.895 207.485 99.045 207.655 ;
        RECT 62.895 204.635 63.425 207.485 ;
        RECT 64.155 206.795 80.155 206.965 ;
        RECT 63.925 205.540 64.095 206.580 ;
        RECT 80.215 205.540 80.385 206.580 ;
        RECT 64.155 205.155 80.155 205.325 ;
        RECT 80.885 204.635 81.055 207.485 ;
        RECT 81.785 206.795 97.785 206.965 ;
        RECT 81.555 205.540 81.725 206.580 ;
        RECT 97.845 205.540 98.015 206.580 ;
        RECT 81.785 205.155 97.785 205.325 ;
        RECT 98.515 204.635 99.045 207.485 ;
        RECT 62.895 204.465 99.045 204.635 ;
        RECT 62.895 201.615 63.425 204.465 ;
        RECT 64.155 203.775 80.155 203.945 ;
        RECT 63.925 202.520 64.095 203.560 ;
        RECT 80.215 202.520 80.385 203.560 ;
        RECT 64.155 202.135 80.155 202.305 ;
        RECT 80.885 201.615 81.055 204.465 ;
        RECT 81.785 203.775 97.785 203.945 ;
        RECT 81.555 202.520 81.725 203.560 ;
        RECT 97.845 202.520 98.015 203.560 ;
        RECT 81.785 202.135 97.785 202.305 ;
        RECT 98.515 201.615 99.045 204.465 ;
        RECT 62.895 201.445 99.045 201.615 ;
        RECT 62.895 198.595 63.425 201.445 ;
        RECT 64.155 200.755 80.155 200.925 ;
        RECT 63.925 199.500 64.095 200.540 ;
        RECT 80.215 199.500 80.385 200.540 ;
        RECT 64.155 199.115 80.155 199.285 ;
        RECT 80.885 198.595 81.055 201.445 ;
        RECT 81.785 200.755 97.785 200.925 ;
        RECT 81.555 199.500 81.725 200.540 ;
        RECT 97.845 199.500 98.015 200.540 ;
        RECT 81.785 199.115 97.785 199.285 ;
        RECT 98.515 198.595 99.045 201.445 ;
        RECT 62.895 198.425 99.045 198.595 ;
        RECT 62.895 195.575 63.425 198.425 ;
        RECT 64.155 197.735 80.155 197.905 ;
        RECT 63.925 196.480 64.095 197.520 ;
        RECT 80.215 196.480 80.385 197.520 ;
        RECT 64.155 196.095 80.155 196.265 ;
        RECT 80.885 195.575 81.055 198.425 ;
        RECT 81.785 197.735 97.785 197.905 ;
        RECT 81.555 196.480 81.725 197.520 ;
        RECT 97.845 196.480 98.015 197.520 ;
        RECT 81.785 196.095 97.785 196.265 ;
        RECT 98.515 195.575 99.045 198.425 ;
        RECT 62.895 195.405 99.045 195.575 ;
        RECT 62.895 192.555 63.425 195.405 ;
        RECT 64.155 194.715 80.155 194.885 ;
        RECT 63.925 193.460 64.095 194.500 ;
        RECT 80.215 193.460 80.385 194.500 ;
        RECT 64.155 193.075 80.155 193.245 ;
        RECT 80.885 192.555 81.055 195.405 ;
        RECT 81.785 194.715 97.785 194.885 ;
        RECT 81.555 193.460 81.725 194.500 ;
        RECT 97.845 193.460 98.015 194.500 ;
        RECT 81.785 193.075 97.785 193.245 ;
        RECT 98.515 192.555 99.045 195.405 ;
        RECT 62.895 192.385 99.045 192.555 ;
        RECT 62.895 189.535 63.425 192.385 ;
        RECT 64.155 191.695 80.155 191.865 ;
        RECT 63.925 190.440 64.095 191.480 ;
        RECT 80.215 190.440 80.385 191.480 ;
        RECT 64.155 190.055 80.155 190.225 ;
        RECT 80.885 189.535 81.055 192.385 ;
        RECT 81.785 191.695 97.785 191.865 ;
        RECT 81.555 190.440 81.725 191.480 ;
        RECT 97.845 190.440 98.015 191.480 ;
        RECT 81.785 190.055 97.785 190.225 ;
        RECT 98.515 189.535 99.045 192.385 ;
        RECT 62.895 189.365 99.045 189.535 ;
        RECT 16.345 180.680 45.335 180.850 ;
        RECT 62.895 186.515 63.425 189.365 ;
        RECT 64.155 188.675 80.155 188.845 ;
        RECT 63.925 187.420 64.095 188.460 ;
        RECT 80.215 187.420 80.385 188.460 ;
        RECT 64.155 187.035 80.155 187.205 ;
        RECT 80.885 186.515 81.055 189.365 ;
        RECT 81.785 188.675 97.785 188.845 ;
        RECT 81.555 187.420 81.725 188.460 ;
        RECT 97.845 187.420 98.015 188.460 ;
        RECT 81.785 187.035 97.785 187.205 ;
        RECT 98.515 186.515 99.045 189.365 ;
        RECT 62.895 186.345 99.045 186.515 ;
        RECT 62.895 183.495 63.425 186.345 ;
        RECT 64.155 185.655 80.155 185.825 ;
        RECT 63.925 184.400 64.095 185.440 ;
        RECT 80.215 184.400 80.385 185.440 ;
        RECT 64.155 184.015 80.155 184.185 ;
        RECT 80.885 183.495 81.055 186.345 ;
        RECT 81.785 185.655 97.785 185.825 ;
        RECT 81.555 184.400 81.725 185.440 ;
        RECT 97.845 184.400 98.015 185.440 ;
        RECT 81.785 184.015 97.785 184.185 ;
        RECT 98.515 183.495 99.045 186.345 ;
        RECT 62.895 183.325 99.045 183.495 ;
        RECT 62.895 180.475 63.425 183.325 ;
        RECT 64.155 182.635 80.155 182.805 ;
        RECT 63.925 181.380 64.095 182.420 ;
        RECT 80.215 181.380 80.385 182.420 ;
        RECT 64.155 180.995 80.155 181.165 ;
        RECT 80.885 180.475 81.055 183.325 ;
        RECT 81.785 182.635 97.785 182.805 ;
        RECT 81.555 181.380 81.725 182.420 ;
        RECT 97.845 181.380 98.015 182.420 ;
        RECT 81.785 180.995 97.785 181.165 ;
        RECT 98.515 180.475 99.045 183.325 ;
        RECT 102.225 181.020 102.625 222.030 ;
        RECT 108.630 220.425 153.130 220.595 ;
        RECT 108.630 216.575 108.800 220.425 ;
        RECT 109.585 219.735 110.585 219.905 ;
        RECT 110.875 219.735 111.875 219.905 ;
        RECT 109.355 217.480 109.525 219.520 ;
        RECT 110.645 217.480 110.815 219.520 ;
        RECT 111.935 217.480 112.105 219.520 ;
        RECT 109.585 217.095 110.585 217.265 ;
        RECT 110.875 217.095 111.875 217.265 ;
        RECT 112.660 216.575 112.830 220.425 ;
        RECT 113.615 219.735 114.615 219.905 ;
        RECT 114.905 219.735 115.905 219.905 ;
        RECT 113.385 217.480 113.555 219.520 ;
        RECT 114.675 217.480 114.845 219.520 ;
        RECT 115.965 217.480 116.135 219.520 ;
        RECT 113.615 217.095 114.615 217.265 ;
        RECT 114.905 217.095 115.905 217.265 ;
        RECT 116.690 216.575 116.860 220.425 ;
        RECT 117.645 219.735 118.645 219.905 ;
        RECT 118.935 219.735 119.935 219.905 ;
        RECT 117.415 217.480 117.585 219.520 ;
        RECT 118.705 217.480 118.875 219.520 ;
        RECT 119.995 217.480 120.165 219.520 ;
        RECT 117.645 217.095 118.645 217.265 ;
        RECT 118.935 217.095 119.935 217.265 ;
        RECT 120.720 216.575 120.890 220.425 ;
        RECT 121.675 219.735 122.675 219.905 ;
        RECT 122.965 219.735 123.965 219.905 ;
        RECT 121.445 217.480 121.615 219.520 ;
        RECT 122.735 217.480 122.905 219.520 ;
        RECT 124.025 217.480 124.195 219.520 ;
        RECT 121.675 217.095 122.675 217.265 ;
        RECT 122.965 217.095 123.965 217.265 ;
        RECT 124.750 216.575 124.920 220.425 ;
        RECT 125.705 219.735 126.705 219.905 ;
        RECT 126.995 219.735 127.995 219.905 ;
        RECT 125.475 217.480 125.645 219.520 ;
        RECT 126.765 217.480 126.935 219.520 ;
        RECT 128.055 217.480 128.225 219.520 ;
        RECT 125.705 217.095 126.705 217.265 ;
        RECT 126.995 217.095 127.995 217.265 ;
        RECT 128.780 216.575 128.950 220.425 ;
        RECT 129.735 219.735 130.735 219.905 ;
        RECT 131.025 219.735 132.025 219.905 ;
        RECT 129.505 217.480 129.675 219.520 ;
        RECT 130.795 217.480 130.965 219.520 ;
        RECT 132.085 217.480 132.255 219.520 ;
        RECT 129.735 217.095 130.735 217.265 ;
        RECT 131.025 217.095 132.025 217.265 ;
        RECT 132.810 216.575 132.980 220.425 ;
        RECT 133.765 219.735 134.765 219.905 ;
        RECT 135.055 219.735 136.055 219.905 ;
        RECT 133.535 217.480 133.705 219.520 ;
        RECT 134.825 217.480 134.995 219.520 ;
        RECT 136.115 217.480 136.285 219.520 ;
        RECT 133.765 217.095 134.765 217.265 ;
        RECT 135.055 217.095 136.055 217.265 ;
        RECT 136.840 216.575 137.010 220.425 ;
        RECT 137.795 219.735 138.795 219.905 ;
        RECT 139.085 219.735 140.085 219.905 ;
        RECT 137.565 217.480 137.735 219.520 ;
        RECT 138.855 217.480 139.025 219.520 ;
        RECT 140.145 217.480 140.315 219.520 ;
        RECT 137.795 217.095 138.795 217.265 ;
        RECT 139.085 217.095 140.085 217.265 ;
        RECT 140.870 216.575 141.040 220.425 ;
        RECT 141.825 219.735 142.825 219.905 ;
        RECT 143.115 219.735 144.115 219.905 ;
        RECT 141.595 217.480 141.765 219.520 ;
        RECT 142.885 217.480 143.055 219.520 ;
        RECT 144.175 217.480 144.345 219.520 ;
        RECT 141.825 217.095 142.825 217.265 ;
        RECT 143.115 217.095 144.115 217.265 ;
        RECT 144.900 216.575 145.070 220.425 ;
        RECT 145.855 219.735 146.855 219.905 ;
        RECT 147.145 219.735 148.145 219.905 ;
        RECT 145.625 217.480 145.795 219.520 ;
        RECT 146.915 217.480 147.085 219.520 ;
        RECT 148.205 217.480 148.375 219.520 ;
        RECT 145.855 217.095 146.855 217.265 ;
        RECT 147.145 217.095 148.145 217.265 ;
        RECT 148.930 216.575 149.100 220.425 ;
        RECT 149.885 219.735 150.885 219.905 ;
        RECT 151.175 219.735 152.175 219.905 ;
        RECT 149.655 217.480 149.825 219.520 ;
        RECT 150.945 217.480 151.115 219.520 ;
        RECT 152.235 217.480 152.405 219.520 ;
        RECT 149.885 217.095 150.885 217.265 ;
        RECT 151.175 217.095 152.175 217.265 ;
        RECT 152.960 216.575 153.130 220.425 ;
        RECT 108.630 216.405 153.130 216.575 ;
        RECT 108.630 213.455 153.130 213.625 ;
        RECT 108.630 203.605 108.800 213.455 ;
        RECT 109.585 212.765 110.585 212.935 ;
        RECT 110.875 212.765 111.875 212.935 ;
        RECT 109.355 204.510 109.525 212.550 ;
        RECT 110.645 204.510 110.815 212.550 ;
        RECT 111.935 204.510 112.105 212.550 ;
        RECT 109.585 204.125 110.585 204.295 ;
        RECT 110.875 204.125 111.875 204.295 ;
        RECT 112.660 203.605 112.830 213.455 ;
        RECT 113.615 212.765 114.615 212.935 ;
        RECT 114.905 212.765 115.905 212.935 ;
        RECT 113.385 204.510 113.555 212.550 ;
        RECT 114.675 204.510 114.845 212.550 ;
        RECT 115.965 204.510 116.135 212.550 ;
        RECT 113.615 204.125 114.615 204.295 ;
        RECT 114.905 204.125 115.905 204.295 ;
        RECT 116.690 203.605 116.860 213.455 ;
        RECT 117.645 212.765 118.645 212.935 ;
        RECT 118.935 212.765 119.935 212.935 ;
        RECT 117.415 204.510 117.585 212.550 ;
        RECT 118.705 204.510 118.875 212.550 ;
        RECT 119.995 204.510 120.165 212.550 ;
        RECT 117.645 204.125 118.645 204.295 ;
        RECT 118.935 204.125 119.935 204.295 ;
        RECT 120.720 203.605 120.890 213.455 ;
        RECT 121.675 212.765 122.675 212.935 ;
        RECT 122.965 212.765 123.965 212.935 ;
        RECT 121.445 204.510 121.615 212.550 ;
        RECT 122.735 204.510 122.905 212.550 ;
        RECT 124.025 204.510 124.195 212.550 ;
        RECT 121.675 204.125 122.675 204.295 ;
        RECT 122.965 204.125 123.965 204.295 ;
        RECT 124.750 203.605 124.920 213.455 ;
        RECT 125.705 212.765 126.705 212.935 ;
        RECT 126.995 212.765 127.995 212.935 ;
        RECT 125.475 204.510 125.645 212.550 ;
        RECT 126.765 204.510 126.935 212.550 ;
        RECT 128.055 204.510 128.225 212.550 ;
        RECT 125.705 204.125 126.705 204.295 ;
        RECT 126.995 204.125 127.995 204.295 ;
        RECT 128.780 203.605 128.950 213.455 ;
        RECT 129.735 212.765 130.735 212.935 ;
        RECT 131.025 212.765 132.025 212.935 ;
        RECT 129.505 204.510 129.675 212.550 ;
        RECT 130.795 204.510 130.965 212.550 ;
        RECT 132.085 204.510 132.255 212.550 ;
        RECT 129.735 204.125 130.735 204.295 ;
        RECT 131.025 204.125 132.025 204.295 ;
        RECT 132.810 203.605 132.980 213.455 ;
        RECT 133.765 212.765 134.765 212.935 ;
        RECT 135.055 212.765 136.055 212.935 ;
        RECT 133.535 204.510 133.705 212.550 ;
        RECT 134.825 204.510 134.995 212.550 ;
        RECT 136.115 204.510 136.285 212.550 ;
        RECT 133.765 204.125 134.765 204.295 ;
        RECT 135.055 204.125 136.055 204.295 ;
        RECT 136.840 203.605 137.010 213.455 ;
        RECT 137.795 212.765 138.795 212.935 ;
        RECT 139.085 212.765 140.085 212.935 ;
        RECT 137.565 204.510 137.735 212.550 ;
        RECT 138.855 204.510 139.025 212.550 ;
        RECT 140.145 204.510 140.315 212.550 ;
        RECT 137.795 204.125 138.795 204.295 ;
        RECT 139.085 204.125 140.085 204.295 ;
        RECT 140.870 203.605 141.040 213.455 ;
        RECT 141.825 212.765 142.825 212.935 ;
        RECT 143.115 212.765 144.115 212.935 ;
        RECT 141.595 204.510 141.765 212.550 ;
        RECT 142.885 204.510 143.055 212.550 ;
        RECT 144.175 204.510 144.345 212.550 ;
        RECT 141.825 204.125 142.825 204.295 ;
        RECT 143.115 204.125 144.115 204.295 ;
        RECT 144.900 203.605 145.070 213.455 ;
        RECT 145.855 212.765 146.855 212.935 ;
        RECT 147.145 212.765 148.145 212.935 ;
        RECT 145.625 204.510 145.795 212.550 ;
        RECT 146.915 204.510 147.085 212.550 ;
        RECT 148.205 204.510 148.375 212.550 ;
        RECT 145.855 204.125 146.855 204.295 ;
        RECT 147.145 204.125 148.145 204.295 ;
        RECT 148.930 203.605 149.100 213.455 ;
        RECT 149.885 212.765 150.885 212.935 ;
        RECT 151.175 212.765 152.175 212.935 ;
        RECT 149.655 204.510 149.825 212.550 ;
        RECT 150.945 204.510 151.115 212.550 ;
        RECT 152.235 204.510 152.405 212.550 ;
        RECT 149.885 204.125 150.885 204.295 ;
        RECT 151.175 204.125 152.175 204.295 ;
        RECT 152.960 203.605 153.130 213.455 ;
        RECT 108.630 203.435 153.130 203.605 ;
        RECT 165.150 201.405 239.210 201.575 ;
        RECT 108.630 200.740 153.130 200.910 ;
        RECT 108.630 194.980 108.800 200.740 ;
        RECT 109.585 200.050 110.585 200.220 ;
        RECT 110.875 200.050 111.875 200.220 ;
        RECT 109.355 195.840 109.525 199.880 ;
        RECT 110.645 195.840 110.815 199.880 ;
        RECT 111.935 195.840 112.105 199.880 ;
        RECT 109.585 195.500 110.585 195.670 ;
        RECT 110.875 195.500 111.875 195.670 ;
        RECT 112.660 194.980 112.830 200.740 ;
        RECT 113.615 200.050 114.615 200.220 ;
        RECT 114.905 200.050 115.905 200.220 ;
        RECT 113.385 195.840 113.555 199.880 ;
        RECT 114.675 195.840 114.845 199.880 ;
        RECT 115.965 195.840 116.135 199.880 ;
        RECT 113.615 195.500 114.615 195.670 ;
        RECT 114.905 195.500 115.905 195.670 ;
        RECT 116.690 194.980 116.860 200.740 ;
        RECT 117.645 200.050 118.645 200.220 ;
        RECT 118.935 200.050 119.935 200.220 ;
        RECT 117.415 195.840 117.585 199.880 ;
        RECT 118.705 195.840 118.875 199.880 ;
        RECT 119.995 195.840 120.165 199.880 ;
        RECT 117.645 195.500 118.645 195.670 ;
        RECT 118.935 195.500 119.935 195.670 ;
        RECT 120.720 194.980 120.890 200.740 ;
        RECT 121.675 200.050 122.675 200.220 ;
        RECT 122.965 200.050 123.965 200.220 ;
        RECT 121.445 195.840 121.615 199.880 ;
        RECT 122.735 195.840 122.905 199.880 ;
        RECT 124.025 195.840 124.195 199.880 ;
        RECT 121.675 195.500 122.675 195.670 ;
        RECT 122.965 195.500 123.965 195.670 ;
        RECT 124.750 194.980 124.920 200.740 ;
        RECT 125.705 200.050 126.705 200.220 ;
        RECT 126.995 200.050 127.995 200.220 ;
        RECT 125.475 195.840 125.645 199.880 ;
        RECT 126.765 195.840 126.935 199.880 ;
        RECT 128.055 195.840 128.225 199.880 ;
        RECT 125.705 195.500 126.705 195.670 ;
        RECT 126.995 195.500 127.995 195.670 ;
        RECT 128.780 194.980 128.950 200.740 ;
        RECT 129.735 200.050 130.735 200.220 ;
        RECT 131.025 200.050 132.025 200.220 ;
        RECT 129.505 195.840 129.675 199.880 ;
        RECT 130.795 195.840 130.965 199.880 ;
        RECT 132.085 195.840 132.255 199.880 ;
        RECT 129.735 195.500 130.735 195.670 ;
        RECT 131.025 195.500 132.025 195.670 ;
        RECT 132.810 194.980 132.980 200.740 ;
        RECT 133.765 200.050 134.765 200.220 ;
        RECT 135.055 200.050 136.055 200.220 ;
        RECT 133.535 195.840 133.705 199.880 ;
        RECT 134.825 195.840 134.995 199.880 ;
        RECT 136.115 195.840 136.285 199.880 ;
        RECT 133.765 195.500 134.765 195.670 ;
        RECT 135.055 195.500 136.055 195.670 ;
        RECT 136.840 194.980 137.010 200.740 ;
        RECT 137.795 200.050 138.795 200.220 ;
        RECT 139.085 200.050 140.085 200.220 ;
        RECT 137.565 195.840 137.735 199.880 ;
        RECT 138.855 195.840 139.025 199.880 ;
        RECT 140.145 195.840 140.315 199.880 ;
        RECT 137.795 195.500 138.795 195.670 ;
        RECT 139.085 195.500 140.085 195.670 ;
        RECT 140.870 194.980 141.040 200.740 ;
        RECT 141.825 200.050 142.825 200.220 ;
        RECT 143.115 200.050 144.115 200.220 ;
        RECT 141.595 195.840 141.765 199.880 ;
        RECT 142.885 195.840 143.055 199.880 ;
        RECT 144.175 195.840 144.345 199.880 ;
        RECT 141.825 195.500 142.825 195.670 ;
        RECT 143.115 195.500 144.115 195.670 ;
        RECT 144.900 194.980 145.070 200.740 ;
        RECT 145.855 200.050 146.855 200.220 ;
        RECT 147.145 200.050 148.145 200.220 ;
        RECT 145.625 195.840 145.795 199.880 ;
        RECT 146.915 195.840 147.085 199.880 ;
        RECT 148.205 195.840 148.375 199.880 ;
        RECT 145.855 195.500 146.855 195.670 ;
        RECT 147.145 195.500 148.145 195.670 ;
        RECT 148.930 194.980 149.100 200.740 ;
        RECT 149.885 200.050 150.885 200.220 ;
        RECT 151.175 200.050 152.175 200.220 ;
        RECT 149.655 195.840 149.825 199.880 ;
        RECT 150.945 195.840 151.115 199.880 ;
        RECT 152.235 195.840 152.405 199.880 ;
        RECT 149.885 195.500 150.885 195.670 ;
        RECT 151.175 195.500 152.175 195.670 ;
        RECT 152.960 194.980 153.130 200.740 ;
        RECT 165.235 200.315 166.445 201.405 ;
        RECT 165.235 199.605 165.755 200.145 ;
        RECT 165.925 199.775 166.445 200.315 ;
        RECT 166.705 200.475 166.875 201.235 ;
        RECT 167.090 200.645 167.420 201.405 ;
        RECT 166.705 200.305 167.420 200.475 ;
        RECT 167.590 200.330 167.845 201.235 ;
        RECT 166.615 199.755 166.970 200.125 ;
        RECT 167.250 200.095 167.420 200.305 ;
        RECT 167.250 199.765 167.505 200.095 ;
        RECT 165.235 198.855 166.445 199.605 ;
        RECT 167.250 199.575 167.420 199.765 ;
        RECT 167.675 199.600 167.845 200.330 ;
        RECT 168.020 200.255 168.280 201.405 ;
        RECT 168.920 200.255 169.180 201.405 ;
        RECT 169.355 200.330 169.610 201.235 ;
        RECT 169.780 200.645 170.110 201.405 ;
        RECT 170.325 200.475 170.495 201.235 ;
        RECT 170.755 200.970 176.100 201.405 ;
        RECT 166.705 199.405 167.420 199.575 ;
        RECT 166.705 199.025 166.875 199.405 ;
        RECT 167.090 198.855 167.420 199.235 ;
        RECT 167.590 199.025 167.845 199.600 ;
        RECT 168.020 198.855 168.280 199.695 ;
        RECT 168.920 198.855 169.180 199.695 ;
        RECT 169.355 199.600 169.525 200.330 ;
        RECT 169.780 200.305 170.495 200.475 ;
        RECT 169.780 200.095 169.950 200.305 ;
        RECT 169.695 199.765 169.950 200.095 ;
        RECT 169.355 199.025 169.610 199.600 ;
        RECT 169.780 199.575 169.950 199.765 ;
        RECT 170.230 199.755 170.585 200.125 ;
        RECT 169.780 199.405 170.495 199.575 ;
        RECT 169.780 198.855 170.110 199.235 ;
        RECT 170.325 199.025 170.495 199.405 ;
        RECT 172.340 199.400 172.680 200.230 ;
        RECT 174.160 199.720 174.510 200.970 ;
        RECT 176.275 200.315 177.945 201.405 ;
        RECT 176.275 199.625 177.025 200.145 ;
        RECT 177.195 199.795 177.945 200.315 ;
        RECT 178.115 200.240 178.405 201.405 ;
        RECT 178.665 200.475 178.835 201.235 ;
        RECT 179.050 200.645 179.380 201.405 ;
        RECT 178.665 200.305 179.380 200.475 ;
        RECT 179.550 200.330 179.805 201.235 ;
        RECT 178.575 199.755 178.930 200.125 ;
        RECT 179.210 200.095 179.380 200.305 ;
        RECT 179.210 199.765 179.465 200.095 ;
        RECT 170.755 198.855 176.100 199.400 ;
        RECT 176.275 198.855 177.945 199.625 ;
        RECT 178.115 198.855 178.405 199.580 ;
        RECT 179.210 199.575 179.380 199.765 ;
        RECT 179.635 199.600 179.805 200.330 ;
        RECT 179.980 200.255 180.240 201.405 ;
        RECT 180.415 200.970 185.760 201.405 ;
        RECT 178.665 199.405 179.380 199.575 ;
        RECT 178.665 199.025 178.835 199.405 ;
        RECT 179.050 198.855 179.380 199.235 ;
        RECT 179.550 199.025 179.805 199.600 ;
        RECT 179.980 198.855 180.240 199.695 ;
        RECT 182.000 199.400 182.340 200.230 ;
        RECT 183.820 199.720 184.170 200.970 ;
        RECT 185.935 200.315 187.605 201.405 ;
        RECT 185.935 199.625 186.685 200.145 ;
        RECT 186.855 199.795 187.605 200.315 ;
        RECT 188.240 200.255 188.500 201.405 ;
        RECT 188.675 200.330 188.930 201.235 ;
        RECT 189.100 200.645 189.430 201.405 ;
        RECT 189.645 200.475 189.815 201.235 ;
        RECT 180.415 198.855 185.760 199.400 ;
        RECT 185.935 198.855 187.605 199.625 ;
        RECT 188.240 198.855 188.500 199.695 ;
        RECT 188.675 199.600 188.845 200.330 ;
        RECT 189.100 200.305 189.815 200.475 ;
        RECT 189.100 200.095 189.270 200.305 ;
        RECT 190.995 200.240 191.285 201.405 ;
        RECT 191.455 200.970 196.800 201.405 ;
        RECT 189.015 199.765 189.270 200.095 ;
        RECT 188.675 199.025 188.930 199.600 ;
        RECT 189.100 199.575 189.270 199.765 ;
        RECT 189.550 199.755 189.905 200.125 ;
        RECT 189.100 199.405 189.815 199.575 ;
        RECT 189.100 198.855 189.430 199.235 ;
        RECT 189.645 199.025 189.815 199.405 ;
        RECT 190.995 198.855 191.285 199.580 ;
        RECT 193.040 199.400 193.380 200.230 ;
        RECT 194.860 199.720 195.210 200.970 ;
        RECT 197.985 200.475 198.155 201.235 ;
        RECT 198.370 200.645 198.700 201.405 ;
        RECT 197.985 200.305 198.700 200.475 ;
        RECT 198.870 200.330 199.125 201.235 ;
        RECT 197.895 199.755 198.250 200.125 ;
        RECT 198.530 200.095 198.700 200.305 ;
        RECT 198.530 199.765 198.785 200.095 ;
        RECT 198.530 199.575 198.700 199.765 ;
        RECT 198.955 199.600 199.125 200.330 ;
        RECT 199.300 200.255 199.560 201.405 ;
        RECT 199.735 200.315 203.245 201.405 ;
        RECT 197.985 199.405 198.700 199.575 ;
        RECT 191.455 198.855 196.800 199.400 ;
        RECT 197.985 199.025 198.155 199.405 ;
        RECT 198.370 198.855 198.700 199.235 ;
        RECT 198.870 199.025 199.125 199.600 ;
        RECT 199.300 198.855 199.560 199.695 ;
        RECT 199.735 199.625 201.385 200.145 ;
        RECT 201.555 199.795 203.245 200.315 ;
        RECT 203.875 200.240 204.165 201.405 ;
        RECT 204.335 200.315 206.925 201.405 ;
        RECT 204.335 199.625 205.545 200.145 ;
        RECT 205.715 199.795 206.925 200.315 ;
        RECT 207.560 200.255 207.820 201.405 ;
        RECT 207.995 200.330 208.250 201.235 ;
        RECT 208.420 200.645 208.750 201.405 ;
        RECT 208.965 200.475 209.135 201.235 ;
        RECT 209.395 200.970 214.740 201.405 ;
        RECT 199.735 198.855 203.245 199.625 ;
        RECT 203.875 198.855 204.165 199.580 ;
        RECT 204.335 198.855 206.925 199.625 ;
        RECT 207.560 198.855 207.820 199.695 ;
        RECT 207.995 199.600 208.165 200.330 ;
        RECT 208.420 200.305 209.135 200.475 ;
        RECT 208.420 200.095 208.590 200.305 ;
        RECT 208.335 199.765 208.590 200.095 ;
        RECT 207.995 199.025 208.250 199.600 ;
        RECT 208.420 199.575 208.590 199.765 ;
        RECT 208.870 199.755 209.225 200.125 ;
        RECT 208.420 199.405 209.135 199.575 ;
        RECT 208.420 198.855 208.750 199.235 ;
        RECT 208.965 199.025 209.135 199.405 ;
        RECT 210.980 199.400 211.320 200.230 ;
        RECT 212.800 199.720 213.150 200.970 ;
        RECT 214.915 200.315 216.585 201.405 ;
        RECT 214.915 199.625 215.665 200.145 ;
        RECT 215.835 199.795 216.585 200.315 ;
        RECT 216.755 200.240 217.045 201.405 ;
        RECT 217.305 200.475 217.475 201.235 ;
        RECT 217.690 200.645 218.020 201.405 ;
        RECT 217.305 200.305 218.020 200.475 ;
        RECT 218.190 200.330 218.445 201.235 ;
        RECT 217.215 199.755 217.570 200.125 ;
        RECT 217.850 200.095 218.020 200.305 ;
        RECT 217.850 199.765 218.105 200.095 ;
        RECT 209.395 198.855 214.740 199.400 ;
        RECT 214.915 198.855 216.585 199.625 ;
        RECT 216.755 198.855 217.045 199.580 ;
        RECT 217.850 199.575 218.020 199.765 ;
        RECT 218.275 199.600 218.445 200.330 ;
        RECT 218.620 200.255 218.880 201.405 ;
        RECT 219.055 200.970 224.400 201.405 ;
        RECT 217.305 199.405 218.020 199.575 ;
        RECT 217.305 199.025 217.475 199.405 ;
        RECT 217.690 198.855 218.020 199.235 ;
        RECT 218.190 199.025 218.445 199.600 ;
        RECT 218.620 198.855 218.880 199.695 ;
        RECT 220.640 199.400 220.980 200.230 ;
        RECT 222.460 199.720 222.810 200.970 ;
        RECT 224.575 200.315 226.245 201.405 ;
        RECT 224.575 199.625 225.325 200.145 ;
        RECT 225.495 199.795 226.245 200.315 ;
        RECT 226.965 200.475 227.135 201.235 ;
        RECT 227.350 200.645 227.680 201.405 ;
        RECT 226.965 200.305 227.680 200.475 ;
        RECT 227.850 200.330 228.105 201.235 ;
        RECT 226.875 199.755 227.230 200.125 ;
        RECT 227.510 200.095 227.680 200.305 ;
        RECT 227.510 199.765 227.765 200.095 ;
        RECT 219.055 198.855 224.400 199.400 ;
        RECT 224.575 198.855 226.245 199.625 ;
        RECT 227.510 199.575 227.680 199.765 ;
        RECT 227.935 199.600 228.105 200.330 ;
        RECT 228.280 200.255 228.540 201.405 ;
        RECT 229.635 200.240 229.925 201.405 ;
        RECT 230.095 200.970 235.440 201.405 ;
        RECT 226.965 199.405 227.680 199.575 ;
        RECT 226.965 199.025 227.135 199.405 ;
        RECT 227.350 198.855 227.680 199.235 ;
        RECT 227.850 199.025 228.105 199.600 ;
        RECT 228.280 198.855 228.540 199.695 ;
        RECT 229.635 198.855 229.925 199.580 ;
        RECT 231.680 199.400 232.020 200.230 ;
        RECT 233.500 199.720 233.850 200.970 ;
        RECT 236.165 200.475 236.335 201.235 ;
        RECT 236.550 200.645 236.880 201.405 ;
        RECT 236.165 200.305 236.880 200.475 ;
        RECT 237.050 200.330 237.305 201.235 ;
        RECT 236.075 199.755 236.430 200.125 ;
        RECT 236.710 200.095 236.880 200.305 ;
        RECT 236.710 199.765 236.965 200.095 ;
        RECT 236.710 199.575 236.880 199.765 ;
        RECT 237.135 199.600 237.305 200.330 ;
        RECT 237.480 200.255 237.740 201.405 ;
        RECT 237.915 200.315 239.125 201.405 ;
        RECT 237.915 199.775 238.435 200.315 ;
        RECT 236.165 199.405 236.880 199.575 ;
        RECT 230.095 198.855 235.440 199.400 ;
        RECT 236.165 199.025 236.335 199.405 ;
        RECT 236.550 198.855 236.880 199.235 ;
        RECT 237.050 199.025 237.305 199.600 ;
        RECT 237.480 198.855 237.740 199.695 ;
        RECT 238.605 199.605 239.125 200.145 ;
        RECT 237.915 198.855 239.125 199.605 ;
        RECT 165.150 198.685 239.210 198.855 ;
        RECT 165.235 197.935 166.445 198.685 ;
        RECT 166.615 198.140 171.960 198.685 ;
        RECT 172.135 198.140 177.480 198.685 ;
        RECT 177.655 198.140 183.000 198.685 ;
        RECT 183.175 198.140 188.520 198.685 ;
        RECT 165.235 197.395 165.755 197.935 ;
        RECT 165.925 197.225 166.445 197.765 ;
        RECT 168.200 197.310 168.540 198.140 ;
        RECT 165.235 196.135 166.445 197.225 ;
        RECT 170.020 196.570 170.370 197.820 ;
        RECT 173.720 197.310 174.060 198.140 ;
        RECT 175.540 196.570 175.890 197.820 ;
        RECT 179.240 197.310 179.580 198.140 ;
        RECT 181.060 196.570 181.410 197.820 ;
        RECT 184.760 197.310 185.100 198.140 ;
        RECT 188.695 197.915 190.365 198.685 ;
        RECT 190.995 197.960 191.285 198.685 ;
        RECT 191.455 198.140 196.800 198.685 ;
        RECT 196.975 198.140 202.320 198.685 ;
        RECT 202.495 198.140 207.840 198.685 ;
        RECT 208.015 198.140 213.360 198.685 ;
        RECT 186.580 196.570 186.930 197.820 ;
        RECT 188.695 197.395 189.445 197.915 ;
        RECT 189.615 197.225 190.365 197.745 ;
        RECT 193.040 197.310 193.380 198.140 ;
        RECT 166.615 196.135 171.960 196.570 ;
        RECT 172.135 196.135 177.480 196.570 ;
        RECT 177.655 196.135 183.000 196.570 ;
        RECT 183.175 196.135 188.520 196.570 ;
        RECT 188.695 196.135 190.365 197.225 ;
        RECT 190.995 196.135 191.285 197.300 ;
        RECT 194.860 196.570 195.210 197.820 ;
        RECT 198.560 197.310 198.900 198.140 ;
        RECT 200.380 196.570 200.730 197.820 ;
        RECT 204.080 197.310 204.420 198.140 ;
        RECT 205.900 196.570 206.250 197.820 ;
        RECT 209.600 197.310 209.940 198.140 ;
        RECT 213.535 197.915 216.125 198.685 ;
        RECT 216.755 197.960 217.045 198.685 ;
        RECT 217.215 198.140 222.560 198.685 ;
        RECT 222.735 198.140 228.080 198.685 ;
        RECT 228.255 198.140 233.600 198.685 ;
        RECT 211.420 196.570 211.770 197.820 ;
        RECT 213.535 197.395 214.745 197.915 ;
        RECT 214.915 197.225 216.125 197.745 ;
        RECT 218.800 197.310 219.140 198.140 ;
        RECT 191.455 196.135 196.800 196.570 ;
        RECT 196.975 196.135 202.320 196.570 ;
        RECT 202.495 196.135 207.840 196.570 ;
        RECT 208.015 196.135 213.360 196.570 ;
        RECT 213.535 196.135 216.125 197.225 ;
        RECT 216.755 196.135 217.045 197.300 ;
        RECT 220.620 196.570 220.970 197.820 ;
        RECT 224.320 197.310 224.660 198.140 ;
        RECT 226.140 196.570 226.490 197.820 ;
        RECT 229.840 197.310 230.180 198.140 ;
        RECT 233.775 197.915 237.285 198.685 ;
        RECT 237.915 197.935 239.125 198.685 ;
        RECT 231.660 196.570 232.010 197.820 ;
        RECT 233.775 197.395 235.425 197.915 ;
        RECT 235.595 197.225 237.285 197.745 ;
        RECT 217.215 196.135 222.560 196.570 ;
        RECT 222.735 196.135 228.080 196.570 ;
        RECT 228.255 196.135 233.600 196.570 ;
        RECT 233.775 196.135 237.285 197.225 ;
        RECT 237.915 197.225 238.435 197.765 ;
        RECT 238.605 197.395 239.125 197.935 ;
        RECT 237.915 196.135 239.125 197.225 ;
        RECT 165.150 195.965 239.210 196.135 ;
        RECT 108.630 194.810 153.130 194.980 ;
        RECT 165.235 194.875 166.445 195.965 ;
        RECT 166.615 195.530 171.960 195.965 ;
        RECT 172.135 195.530 177.480 195.965 ;
        RECT 108.630 185.050 108.800 194.810 ;
        RECT 109.585 194.120 110.585 194.290 ;
        RECT 110.875 194.120 111.875 194.290 ;
        RECT 109.355 185.910 109.525 193.950 ;
        RECT 110.645 185.910 110.815 193.950 ;
        RECT 111.935 185.910 112.105 193.950 ;
        RECT 109.585 185.570 110.585 185.740 ;
        RECT 110.875 185.570 111.875 185.740 ;
        RECT 112.660 185.050 112.830 194.810 ;
        RECT 113.615 194.120 114.615 194.290 ;
        RECT 114.905 194.120 115.905 194.290 ;
        RECT 113.385 185.910 113.555 193.950 ;
        RECT 114.675 185.910 114.845 193.950 ;
        RECT 115.965 185.910 116.135 193.950 ;
        RECT 113.615 185.570 114.615 185.740 ;
        RECT 114.905 185.570 115.905 185.740 ;
        RECT 116.690 185.050 116.860 194.810 ;
        RECT 117.645 194.120 118.645 194.290 ;
        RECT 118.935 194.120 119.935 194.290 ;
        RECT 117.415 185.910 117.585 193.950 ;
        RECT 118.705 185.910 118.875 193.950 ;
        RECT 119.995 185.910 120.165 193.950 ;
        RECT 117.645 185.570 118.645 185.740 ;
        RECT 118.935 185.570 119.935 185.740 ;
        RECT 120.720 185.050 120.890 194.810 ;
        RECT 121.675 194.120 122.675 194.290 ;
        RECT 122.965 194.120 123.965 194.290 ;
        RECT 121.445 185.910 121.615 193.950 ;
        RECT 122.735 185.910 122.905 193.950 ;
        RECT 124.025 185.910 124.195 193.950 ;
        RECT 121.675 185.570 122.675 185.740 ;
        RECT 122.965 185.570 123.965 185.740 ;
        RECT 124.750 185.050 124.920 194.810 ;
        RECT 125.705 194.120 126.705 194.290 ;
        RECT 126.995 194.120 127.995 194.290 ;
        RECT 125.475 185.910 125.645 193.950 ;
        RECT 126.765 185.910 126.935 193.950 ;
        RECT 128.055 185.910 128.225 193.950 ;
        RECT 125.705 185.570 126.705 185.740 ;
        RECT 126.995 185.570 127.995 185.740 ;
        RECT 128.780 185.050 128.950 194.810 ;
        RECT 129.735 194.120 130.735 194.290 ;
        RECT 131.025 194.120 132.025 194.290 ;
        RECT 129.505 185.910 129.675 193.950 ;
        RECT 130.795 185.910 130.965 193.950 ;
        RECT 132.085 185.910 132.255 193.950 ;
        RECT 129.735 185.570 130.735 185.740 ;
        RECT 131.025 185.570 132.025 185.740 ;
        RECT 132.810 185.050 132.980 194.810 ;
        RECT 133.765 194.120 134.765 194.290 ;
        RECT 135.055 194.120 136.055 194.290 ;
        RECT 133.535 185.910 133.705 193.950 ;
        RECT 134.825 185.910 134.995 193.950 ;
        RECT 136.115 185.910 136.285 193.950 ;
        RECT 133.765 185.570 134.765 185.740 ;
        RECT 135.055 185.570 136.055 185.740 ;
        RECT 136.840 185.050 137.010 194.810 ;
        RECT 137.795 194.120 138.795 194.290 ;
        RECT 139.085 194.120 140.085 194.290 ;
        RECT 137.565 185.910 137.735 193.950 ;
        RECT 138.855 185.910 139.025 193.950 ;
        RECT 140.145 185.910 140.315 193.950 ;
        RECT 137.795 185.570 138.795 185.740 ;
        RECT 139.085 185.570 140.085 185.740 ;
        RECT 140.870 185.050 141.040 194.810 ;
        RECT 141.825 194.120 142.825 194.290 ;
        RECT 143.115 194.120 144.115 194.290 ;
        RECT 141.595 185.910 141.765 193.950 ;
        RECT 142.885 185.910 143.055 193.950 ;
        RECT 144.175 185.910 144.345 193.950 ;
        RECT 141.825 185.570 142.825 185.740 ;
        RECT 143.115 185.570 144.115 185.740 ;
        RECT 144.900 185.050 145.070 194.810 ;
        RECT 145.855 194.120 146.855 194.290 ;
        RECT 147.145 194.120 148.145 194.290 ;
        RECT 145.625 185.910 145.795 193.950 ;
        RECT 146.915 185.910 147.085 193.950 ;
        RECT 148.205 185.910 148.375 193.950 ;
        RECT 145.855 185.570 146.855 185.740 ;
        RECT 147.145 185.570 148.145 185.740 ;
        RECT 148.930 185.050 149.100 194.810 ;
        RECT 149.885 194.120 150.885 194.290 ;
        RECT 151.175 194.120 152.175 194.290 ;
        RECT 149.655 185.910 149.825 193.950 ;
        RECT 150.945 185.910 151.115 193.950 ;
        RECT 152.235 185.910 152.405 193.950 ;
        RECT 149.885 185.570 150.885 185.740 ;
        RECT 151.175 185.570 152.175 185.740 ;
        RECT 152.960 185.050 153.130 194.810 ;
        RECT 165.235 194.165 165.755 194.705 ;
        RECT 165.925 194.335 166.445 194.875 ;
        RECT 165.235 193.415 166.445 194.165 ;
        RECT 168.200 193.960 168.540 194.790 ;
        RECT 170.020 194.280 170.370 195.530 ;
        RECT 173.720 193.960 174.060 194.790 ;
        RECT 175.540 194.280 175.890 195.530 ;
        RECT 178.115 194.800 178.405 195.965 ;
        RECT 178.575 195.530 183.920 195.965 ;
        RECT 184.095 195.530 189.440 195.965 ;
        RECT 189.615 195.530 194.960 195.965 ;
        RECT 195.135 195.530 200.480 195.965 ;
        RECT 166.615 193.415 171.960 193.960 ;
        RECT 172.135 193.415 177.480 193.960 ;
        RECT 178.115 193.415 178.405 194.140 ;
        RECT 180.160 193.960 180.500 194.790 ;
        RECT 181.980 194.280 182.330 195.530 ;
        RECT 185.680 193.960 186.020 194.790 ;
        RECT 187.500 194.280 187.850 195.530 ;
        RECT 191.200 193.960 191.540 194.790 ;
        RECT 193.020 194.280 193.370 195.530 ;
        RECT 196.720 193.960 197.060 194.790 ;
        RECT 198.540 194.280 198.890 195.530 ;
        RECT 200.655 194.875 203.245 195.965 ;
        RECT 200.655 194.185 201.865 194.705 ;
        RECT 202.035 194.355 203.245 194.875 ;
        RECT 203.875 194.800 204.165 195.965 ;
        RECT 204.335 195.530 209.680 195.965 ;
        RECT 209.855 195.530 215.200 195.965 ;
        RECT 215.375 195.530 220.720 195.965 ;
        RECT 220.895 195.530 226.240 195.965 ;
        RECT 178.575 193.415 183.920 193.960 ;
        RECT 184.095 193.415 189.440 193.960 ;
        RECT 189.615 193.415 194.960 193.960 ;
        RECT 195.135 193.415 200.480 193.960 ;
        RECT 200.655 193.415 203.245 194.185 ;
        RECT 203.875 193.415 204.165 194.140 ;
        RECT 205.920 193.960 206.260 194.790 ;
        RECT 207.740 194.280 208.090 195.530 ;
        RECT 211.440 193.960 211.780 194.790 ;
        RECT 213.260 194.280 213.610 195.530 ;
        RECT 216.960 193.960 217.300 194.790 ;
        RECT 218.780 194.280 219.130 195.530 ;
        RECT 222.480 193.960 222.820 194.790 ;
        RECT 224.300 194.280 224.650 195.530 ;
        RECT 226.415 194.875 229.005 195.965 ;
        RECT 226.415 194.185 227.625 194.705 ;
        RECT 227.795 194.355 229.005 194.875 ;
        RECT 229.635 194.800 229.925 195.965 ;
        RECT 230.095 195.530 235.440 195.965 ;
        RECT 204.335 193.415 209.680 193.960 ;
        RECT 209.855 193.415 215.200 193.960 ;
        RECT 215.375 193.415 220.720 193.960 ;
        RECT 220.895 193.415 226.240 193.960 ;
        RECT 226.415 193.415 229.005 194.185 ;
        RECT 229.635 193.415 229.925 194.140 ;
        RECT 231.680 193.960 232.020 194.790 ;
        RECT 233.500 194.280 233.850 195.530 ;
        RECT 235.615 194.875 237.285 195.965 ;
        RECT 235.615 194.185 236.365 194.705 ;
        RECT 236.535 194.355 237.285 194.875 ;
        RECT 237.915 194.875 239.125 195.965 ;
        RECT 237.915 194.335 238.435 194.875 ;
        RECT 230.095 193.415 235.440 193.960 ;
        RECT 235.615 193.415 237.285 194.185 ;
        RECT 238.605 194.165 239.125 194.705 ;
        RECT 237.915 193.415 239.125 194.165 ;
        RECT 165.150 193.245 239.210 193.415 ;
        RECT 165.235 192.495 166.445 193.245 ;
        RECT 166.615 192.700 171.960 193.245 ;
        RECT 165.235 191.955 165.755 192.495 ;
        RECT 165.925 191.785 166.445 192.325 ;
        RECT 168.200 191.870 168.540 192.700 ;
        RECT 173.055 192.570 173.315 193.075 ;
        RECT 173.495 192.865 173.825 193.245 ;
        RECT 174.005 192.695 174.175 193.075 ;
        RECT 165.235 190.695 166.445 191.785 ;
        RECT 170.020 191.130 170.370 192.380 ;
        RECT 173.055 191.770 173.225 192.570 ;
        RECT 173.510 192.525 174.175 192.695 ;
        RECT 174.525 192.695 174.695 193.075 ;
        RECT 174.875 192.865 175.205 193.245 ;
        RECT 174.525 192.525 175.190 192.695 ;
        RECT 175.385 192.570 175.645 193.075 ;
        RECT 175.820 192.845 176.155 193.245 ;
        RECT 176.325 192.675 176.530 193.075 ;
        RECT 176.740 192.765 177.015 193.245 ;
        RECT 177.225 192.745 177.485 193.075 ;
        RECT 173.510 192.270 173.680 192.525 ;
        RECT 173.395 191.940 173.680 192.270 ;
        RECT 173.915 191.975 174.245 192.345 ;
        RECT 174.455 191.975 174.785 192.345 ;
        RECT 175.020 192.270 175.190 192.525 ;
        RECT 173.510 191.795 173.680 191.940 ;
        RECT 175.020 191.940 175.305 192.270 ;
        RECT 175.020 191.795 175.190 191.940 ;
        RECT 166.615 190.695 171.960 191.130 ;
        RECT 173.055 190.865 173.325 191.770 ;
        RECT 173.510 191.625 174.175 191.795 ;
        RECT 173.495 190.695 173.825 191.455 ;
        RECT 174.005 190.865 174.175 191.625 ;
        RECT 174.525 191.625 175.190 191.795 ;
        RECT 175.475 191.770 175.645 192.570 ;
        RECT 174.525 190.865 174.695 191.625 ;
        RECT 174.875 190.695 175.205 191.455 ;
        RECT 175.375 190.865 175.645 191.770 ;
        RECT 175.845 192.505 176.530 192.675 ;
        RECT 175.845 191.475 176.185 192.505 ;
        RECT 176.355 191.835 176.605 192.335 ;
        RECT 176.785 192.005 177.145 192.585 ;
        RECT 177.315 191.835 177.485 192.745 ;
        RECT 176.355 191.665 177.485 191.835 ;
        RECT 175.845 191.300 176.510 191.475 ;
        RECT 175.820 190.695 176.155 191.120 ;
        RECT 176.325 190.895 176.510 191.300 ;
        RECT 176.715 190.695 177.045 191.475 ;
        RECT 177.215 190.895 177.485 191.665 ;
        RECT 177.655 192.300 177.995 193.075 ;
        RECT 178.165 192.785 178.335 193.245 ;
        RECT 178.575 192.810 178.935 193.075 ;
        RECT 178.575 192.805 178.930 192.810 ;
        RECT 178.575 192.795 178.925 192.805 ;
        RECT 178.575 192.790 178.920 192.795 ;
        RECT 178.575 192.780 178.915 192.790 ;
        RECT 179.565 192.785 179.735 193.245 ;
        RECT 178.575 192.775 178.910 192.780 ;
        RECT 178.575 192.765 178.900 192.775 ;
        RECT 178.575 192.755 178.890 192.765 ;
        RECT 178.575 192.615 178.875 192.755 ;
        RECT 178.165 192.425 178.875 192.615 ;
        RECT 179.065 192.615 179.395 192.695 ;
        RECT 179.905 192.615 180.245 193.075 ;
        RECT 179.065 192.425 180.245 192.615 ;
        RECT 180.505 192.695 180.675 193.075 ;
        RECT 180.890 192.865 181.220 193.245 ;
        RECT 180.505 192.525 181.220 192.695 ;
        RECT 177.655 190.865 177.935 192.300 ;
        RECT 178.165 191.855 178.450 192.425 ;
        RECT 178.635 192.025 179.105 192.255 ;
        RECT 179.275 192.235 179.605 192.255 ;
        RECT 179.275 192.055 179.725 192.235 ;
        RECT 179.915 192.055 180.245 192.255 ;
        RECT 178.165 191.640 179.315 191.855 ;
        RECT 178.105 190.695 178.815 191.470 ;
        RECT 178.985 190.865 179.315 191.640 ;
        RECT 179.510 190.940 179.725 192.055 ;
        RECT 180.015 191.715 180.245 192.055 ;
        RECT 180.415 191.975 180.770 192.345 ;
        RECT 181.050 192.335 181.220 192.525 ;
        RECT 181.390 192.500 181.645 193.075 ;
        RECT 181.050 192.005 181.305 192.335 ;
        RECT 181.050 191.795 181.220 192.005 ;
        RECT 180.505 191.625 181.220 191.795 ;
        RECT 181.475 191.770 181.645 192.500 ;
        RECT 181.820 192.405 182.080 193.245 ;
        RECT 182.345 192.695 182.515 193.075 ;
        RECT 182.695 192.865 183.025 193.245 ;
        RECT 182.345 192.525 183.010 192.695 ;
        RECT 183.205 192.570 183.465 193.075 ;
        RECT 182.275 191.975 182.605 192.345 ;
        RECT 182.840 192.270 183.010 192.525 ;
        RECT 182.840 191.940 183.125 192.270 ;
        RECT 179.905 190.695 180.235 191.415 ;
        RECT 180.505 190.865 180.675 191.625 ;
        RECT 180.890 190.695 181.220 191.455 ;
        RECT 181.390 190.865 181.645 191.770 ;
        RECT 181.820 190.695 182.080 191.845 ;
        RECT 182.840 191.795 183.010 191.940 ;
        RECT 182.345 191.625 183.010 191.795 ;
        RECT 183.295 191.770 183.465 192.570 ;
        RECT 184.185 192.595 184.355 193.075 ;
        RECT 184.525 192.765 184.855 193.245 ;
        RECT 185.080 192.825 186.615 193.075 ;
        RECT 185.080 192.595 185.250 192.825 ;
        RECT 184.185 192.425 185.250 192.595 ;
        RECT 185.430 192.255 185.710 192.655 ;
        RECT 184.100 192.045 184.450 192.255 ;
        RECT 184.620 192.055 185.065 192.255 ;
        RECT 185.235 192.055 185.710 192.255 ;
        RECT 185.980 192.255 186.265 192.655 ;
        RECT 186.445 192.595 186.615 192.825 ;
        RECT 186.785 192.765 187.115 193.245 ;
        RECT 187.330 192.745 187.585 193.075 ;
        RECT 187.400 192.665 187.585 192.745 ;
        RECT 186.445 192.425 187.245 192.595 ;
        RECT 185.980 192.055 186.310 192.255 ;
        RECT 186.480 192.055 186.845 192.255 ;
        RECT 187.075 191.875 187.245 192.425 ;
        RECT 182.345 190.865 182.515 191.625 ;
        RECT 182.695 190.695 183.025 191.455 ;
        RECT 183.195 190.865 183.465 191.770 ;
        RECT 184.185 191.705 187.245 191.875 ;
        RECT 184.185 190.865 184.355 191.705 ;
        RECT 187.415 191.545 187.585 192.665 ;
        RECT 187.775 192.475 190.365 193.245 ;
        RECT 190.995 192.520 191.285 193.245 ;
        RECT 187.775 191.955 188.985 192.475 ;
        RECT 189.155 191.785 190.365 192.305 ;
        RECT 191.455 192.300 191.795 193.075 ;
        RECT 191.965 192.785 192.135 193.245 ;
        RECT 192.375 192.810 192.735 193.075 ;
        RECT 192.375 192.805 192.730 192.810 ;
        RECT 192.375 192.795 192.725 192.805 ;
        RECT 192.375 192.790 192.720 192.795 ;
        RECT 192.375 192.780 192.715 192.790 ;
        RECT 193.365 192.785 193.535 193.245 ;
        RECT 192.375 192.775 192.710 192.780 ;
        RECT 192.375 192.765 192.700 192.775 ;
        RECT 192.375 192.755 192.690 192.765 ;
        RECT 192.375 192.615 192.675 192.755 ;
        RECT 191.965 192.425 192.675 192.615 ;
        RECT 192.865 192.615 193.195 192.695 ;
        RECT 193.705 192.615 194.045 193.075 ;
        RECT 192.865 192.425 194.045 192.615 ;
        RECT 194.215 192.475 195.885 193.245 ;
        RECT 187.375 191.535 187.585 191.545 ;
        RECT 184.525 191.035 184.855 191.535 ;
        RECT 185.025 191.295 186.660 191.535 ;
        RECT 185.025 191.205 185.255 191.295 ;
        RECT 185.365 191.035 185.695 191.075 ;
        RECT 184.525 190.865 185.695 191.035 ;
        RECT 185.885 190.695 186.240 191.115 ;
        RECT 186.410 190.865 186.660 191.295 ;
        RECT 186.830 190.695 187.160 191.455 ;
        RECT 187.330 190.865 187.585 191.535 ;
        RECT 187.775 190.695 190.365 191.785 ;
        RECT 190.995 190.695 191.285 191.860 ;
        RECT 191.455 190.865 191.735 192.300 ;
        RECT 191.965 191.855 192.250 192.425 ;
        RECT 192.435 192.025 192.905 192.255 ;
        RECT 193.075 192.235 193.405 192.255 ;
        RECT 193.075 192.055 193.525 192.235 ;
        RECT 193.715 192.055 194.045 192.255 ;
        RECT 191.965 191.640 193.115 191.855 ;
        RECT 191.905 190.695 192.615 191.470 ;
        RECT 192.785 190.865 193.115 191.640 ;
        RECT 193.310 190.940 193.525 192.055 ;
        RECT 193.815 191.715 194.045 192.055 ;
        RECT 194.215 191.955 194.965 192.475 ;
        RECT 196.575 192.425 196.785 193.245 ;
        RECT 196.955 192.445 197.285 193.075 ;
        RECT 195.135 191.785 195.885 192.305 ;
        RECT 196.955 191.845 197.205 192.445 ;
        RECT 197.455 192.425 197.685 193.245 ;
        RECT 197.895 192.300 198.235 193.075 ;
        RECT 198.405 192.785 198.575 193.245 ;
        RECT 198.815 192.810 199.175 193.075 ;
        RECT 198.815 192.805 199.170 192.810 ;
        RECT 198.815 192.795 199.165 192.805 ;
        RECT 198.815 192.790 199.160 192.795 ;
        RECT 198.815 192.780 199.155 192.790 ;
        RECT 199.805 192.785 199.975 193.245 ;
        RECT 198.815 192.775 199.150 192.780 ;
        RECT 198.815 192.765 199.140 192.775 ;
        RECT 198.815 192.755 199.130 192.765 ;
        RECT 198.815 192.615 199.115 192.755 ;
        RECT 198.405 192.425 199.115 192.615 ;
        RECT 199.305 192.615 199.635 192.695 ;
        RECT 200.145 192.615 200.485 193.075 ;
        RECT 200.655 192.700 206.000 193.245 ;
        RECT 206.175 192.700 211.520 193.245 ;
        RECT 199.305 192.425 200.485 192.615 ;
        RECT 197.375 192.005 197.705 192.255 ;
        RECT 193.705 190.695 194.035 191.415 ;
        RECT 194.215 190.695 195.885 191.785 ;
        RECT 196.575 190.695 196.785 191.835 ;
        RECT 196.955 190.865 197.285 191.845 ;
        RECT 197.455 190.695 197.685 191.835 ;
        RECT 197.895 190.865 198.175 192.300 ;
        RECT 198.405 191.855 198.690 192.425 ;
        RECT 198.875 192.025 199.345 192.255 ;
        RECT 199.515 192.235 199.845 192.255 ;
        RECT 199.515 192.055 199.965 192.235 ;
        RECT 200.155 192.055 200.485 192.255 ;
        RECT 198.405 191.640 199.555 191.855 ;
        RECT 198.345 190.695 199.055 191.470 ;
        RECT 199.225 190.865 199.555 191.640 ;
        RECT 199.750 190.940 199.965 192.055 ;
        RECT 200.255 191.715 200.485 192.055 ;
        RECT 202.240 191.870 202.580 192.700 ;
        RECT 200.145 190.695 200.475 191.415 ;
        RECT 204.060 191.130 204.410 192.380 ;
        RECT 207.760 191.870 208.100 192.700 ;
        RECT 211.695 192.475 215.205 193.245 ;
        RECT 215.375 192.495 216.585 193.245 ;
        RECT 216.755 192.520 217.045 193.245 ;
        RECT 217.215 192.700 222.560 193.245 ;
        RECT 222.735 192.700 228.080 193.245 ;
        RECT 228.255 192.700 233.600 193.245 ;
        RECT 209.580 191.130 209.930 192.380 ;
        RECT 211.695 191.955 213.345 192.475 ;
        RECT 213.515 191.785 215.205 192.305 ;
        RECT 215.375 191.955 215.895 192.495 ;
        RECT 216.065 191.785 216.585 192.325 ;
        RECT 218.800 191.870 219.140 192.700 ;
        RECT 200.655 190.695 206.000 191.130 ;
        RECT 206.175 190.695 211.520 191.130 ;
        RECT 211.695 190.695 215.205 191.785 ;
        RECT 215.375 190.695 216.585 191.785 ;
        RECT 216.755 190.695 217.045 191.860 ;
        RECT 220.620 191.130 220.970 192.380 ;
        RECT 224.320 191.870 224.660 192.700 ;
        RECT 226.140 191.130 226.490 192.380 ;
        RECT 229.840 191.870 230.180 192.700 ;
        RECT 233.775 192.475 237.285 193.245 ;
        RECT 237.915 192.495 239.125 193.245 ;
        RECT 231.660 191.130 232.010 192.380 ;
        RECT 233.775 191.955 235.425 192.475 ;
        RECT 235.595 191.785 237.285 192.305 ;
        RECT 217.215 190.695 222.560 191.130 ;
        RECT 222.735 190.695 228.080 191.130 ;
        RECT 228.255 190.695 233.600 191.130 ;
        RECT 233.775 190.695 237.285 191.785 ;
        RECT 237.915 191.785 238.435 192.325 ;
        RECT 238.605 191.955 239.125 192.495 ;
        RECT 237.915 190.695 239.125 191.785 ;
        RECT 165.150 190.525 239.210 190.695 ;
        RECT 165.235 189.435 166.445 190.525 ;
        RECT 165.235 188.725 165.755 189.265 ;
        RECT 165.925 188.895 166.445 189.435 ;
        RECT 166.705 189.595 166.875 190.355 ;
        RECT 167.055 189.765 167.385 190.525 ;
        RECT 166.705 189.425 167.370 189.595 ;
        RECT 167.555 189.450 167.825 190.355 ;
        RECT 167.200 189.280 167.370 189.425 ;
        RECT 166.635 188.875 166.965 189.245 ;
        RECT 167.200 188.950 167.485 189.280 ;
        RECT 165.235 187.975 166.445 188.725 ;
        RECT 167.200 188.695 167.370 188.950 ;
        RECT 166.705 188.525 167.370 188.695 ;
        RECT 167.655 188.650 167.825 189.450 ;
        RECT 167.995 189.435 169.665 190.525 ;
        RECT 166.705 188.145 166.875 188.525 ;
        RECT 167.055 187.975 167.385 188.355 ;
        RECT 167.565 188.145 167.825 188.650 ;
        RECT 167.995 188.745 168.745 189.265 ;
        RECT 168.915 188.915 169.665 189.435 ;
        RECT 169.925 189.595 170.095 190.355 ;
        RECT 170.275 189.765 170.605 190.525 ;
        RECT 169.925 189.425 170.590 189.595 ;
        RECT 170.775 189.450 171.045 190.355 ;
        RECT 170.420 189.280 170.590 189.425 ;
        RECT 169.855 188.875 170.185 189.245 ;
        RECT 170.420 188.950 170.705 189.280 ;
        RECT 167.995 187.975 169.665 188.745 ;
        RECT 170.420 188.695 170.590 188.950 ;
        RECT 169.925 188.525 170.590 188.695 ;
        RECT 170.875 188.650 171.045 189.450 ;
        RECT 169.925 188.145 170.095 188.525 ;
        RECT 170.275 187.975 170.605 188.355 ;
        RECT 170.785 188.145 171.045 188.650 ;
        RECT 171.215 188.920 171.495 190.355 ;
        RECT 171.665 189.750 172.375 190.525 ;
        RECT 172.545 189.580 172.875 190.355 ;
        RECT 171.725 189.365 172.875 189.580 ;
        RECT 171.215 188.145 171.555 188.920 ;
        RECT 171.725 188.795 172.010 189.365 ;
        RECT 172.195 188.965 172.665 189.195 ;
        RECT 173.070 189.165 173.285 190.280 ;
        RECT 173.465 189.805 173.795 190.525 ;
        RECT 173.575 189.165 173.805 189.505 ;
        RECT 174.190 189.425 174.520 190.525 ;
        RECT 174.995 189.925 175.320 190.355 ;
        RECT 175.490 190.105 175.820 190.525 ;
        RECT 176.565 190.095 176.975 190.525 ;
        RECT 174.995 189.755 176.975 189.925 ;
        RECT 174.995 189.345 175.700 189.755 ;
        RECT 172.835 188.985 173.285 189.165 ;
        RECT 172.835 188.965 173.165 188.985 ;
        RECT 173.475 188.965 173.805 189.165 ;
        RECT 173.975 188.965 174.620 189.175 ;
        RECT 174.790 188.965 175.360 189.175 ;
        RECT 171.725 188.605 172.435 188.795 ;
        RECT 172.135 188.465 172.435 188.605 ;
        RECT 172.625 188.605 173.805 188.795 ;
        RECT 172.625 188.525 172.955 188.605 ;
        RECT 172.135 188.455 172.450 188.465 ;
        RECT 172.135 188.445 172.460 188.455 ;
        RECT 172.135 188.440 172.470 188.445 ;
        RECT 171.725 187.975 171.895 188.435 ;
        RECT 172.135 188.430 172.475 188.440 ;
        RECT 172.135 188.425 172.480 188.430 ;
        RECT 172.135 188.415 172.485 188.425 ;
        RECT 172.135 188.410 172.490 188.415 ;
        RECT 172.135 188.145 172.495 188.410 ;
        RECT 173.125 187.975 173.295 188.435 ;
        RECT 173.465 188.145 173.805 188.605 ;
        RECT 174.130 188.625 175.300 188.795 ;
        RECT 174.130 188.160 174.460 188.625 ;
        RECT 174.630 187.975 174.800 188.445 ;
        RECT 174.970 188.145 175.300 188.625 ;
        RECT 175.530 188.145 175.700 189.345 ;
        RECT 175.870 189.415 176.495 189.585 ;
        RECT 175.870 188.715 176.040 189.415 ;
        RECT 176.710 189.215 176.975 189.755 ;
        RECT 177.145 189.370 177.485 190.355 ;
        RECT 176.210 188.885 176.540 189.215 ;
        RECT 176.710 188.885 177.060 189.215 ;
        RECT 177.230 188.715 177.485 189.370 ;
        RECT 178.115 189.360 178.405 190.525 ;
        RECT 178.790 189.425 179.120 190.525 ;
        RECT 179.595 189.925 179.920 190.355 ;
        RECT 180.090 190.105 180.420 190.525 ;
        RECT 181.165 190.095 181.575 190.525 ;
        RECT 179.595 189.755 181.575 189.925 ;
        RECT 179.595 189.345 180.300 189.755 ;
        RECT 178.575 188.965 179.220 189.175 ;
        RECT 179.390 188.965 179.960 189.175 ;
        RECT 175.870 188.545 176.410 188.715 ;
        RECT 176.240 188.340 176.410 188.545 ;
        RECT 176.690 187.975 176.860 188.715 ;
        RECT 177.125 188.340 177.485 188.715 ;
        RECT 177.255 188.315 177.425 188.340 ;
        RECT 178.115 187.975 178.405 188.700 ;
        RECT 178.730 188.625 179.900 188.795 ;
        RECT 178.730 188.160 179.060 188.625 ;
        RECT 179.230 187.975 179.400 188.445 ;
        RECT 179.570 188.145 179.900 188.625 ;
        RECT 180.130 188.145 180.300 189.345 ;
        RECT 180.470 189.415 181.095 189.585 ;
        RECT 180.470 188.715 180.640 189.415 ;
        RECT 181.310 189.215 181.575 189.755 ;
        RECT 181.745 189.370 182.085 190.355 ;
        RECT 183.210 189.725 183.460 190.525 ;
        RECT 183.630 189.895 183.960 190.355 ;
        RECT 184.130 190.065 184.345 190.525 ;
        RECT 183.630 189.725 184.800 189.895 ;
        RECT 182.720 189.555 183.000 189.715 ;
        RECT 182.720 189.385 184.055 189.555 ;
        RECT 180.810 188.885 181.140 189.215 ;
        RECT 181.310 188.885 181.660 189.215 ;
        RECT 181.830 188.715 182.085 189.370 ;
        RECT 183.885 189.215 184.055 189.385 ;
        RECT 182.720 188.965 183.070 189.205 ;
        RECT 183.240 188.965 183.715 189.205 ;
        RECT 183.885 188.965 184.260 189.215 ;
        RECT 183.885 188.795 184.055 188.965 ;
        RECT 180.470 188.545 181.010 188.715 ;
        RECT 180.840 188.340 181.010 188.545 ;
        RECT 181.290 187.975 181.460 188.715 ;
        RECT 181.725 188.340 182.085 188.715 ;
        RECT 182.720 188.625 184.055 188.795 ;
        RECT 182.720 188.415 182.990 188.625 ;
        RECT 184.430 188.435 184.800 189.725 ;
        RECT 183.210 187.975 183.540 188.435 ;
        RECT 184.050 188.145 184.800 188.435 ;
        RECT 185.015 189.450 185.285 190.355 ;
        RECT 185.455 189.765 185.785 190.525 ;
        RECT 185.965 189.595 186.135 190.355 ;
        RECT 186.890 189.725 187.140 190.525 ;
        RECT 187.310 189.895 187.640 190.355 ;
        RECT 187.810 190.065 188.025 190.525 ;
        RECT 187.310 189.725 188.480 189.895 ;
        RECT 185.015 188.650 185.185 189.450 ;
        RECT 185.470 189.425 186.135 189.595 ;
        RECT 186.400 189.555 186.680 189.715 ;
        RECT 185.470 189.280 185.640 189.425 ;
        RECT 186.400 189.385 187.735 189.555 ;
        RECT 185.355 188.950 185.640 189.280 ;
        RECT 185.470 188.695 185.640 188.950 ;
        RECT 185.875 188.875 186.205 189.245 ;
        RECT 187.565 189.215 187.735 189.385 ;
        RECT 186.400 188.965 186.750 189.205 ;
        RECT 186.920 188.965 187.395 189.205 ;
        RECT 187.565 188.965 187.940 189.215 ;
        RECT 187.565 188.795 187.735 188.965 ;
        RECT 185.015 188.145 185.275 188.650 ;
        RECT 185.470 188.525 186.135 188.695 ;
        RECT 185.455 187.975 185.785 188.355 ;
        RECT 185.965 188.145 186.135 188.525 ;
        RECT 186.400 188.625 187.735 188.795 ;
        RECT 186.400 188.415 186.670 188.625 ;
        RECT 188.110 188.435 188.480 189.725 ;
        RECT 189.705 189.515 189.875 190.355 ;
        RECT 190.045 190.185 191.215 190.355 ;
        RECT 190.045 189.685 190.375 190.185 ;
        RECT 190.885 190.145 191.215 190.185 ;
        RECT 191.405 190.105 191.760 190.525 ;
        RECT 190.545 189.925 190.775 190.015 ;
        RECT 191.930 189.925 192.180 190.355 ;
        RECT 190.545 189.685 192.180 189.925 ;
        RECT 192.350 189.765 192.680 190.525 ;
        RECT 192.850 189.685 193.105 190.355 ;
        RECT 189.705 189.345 192.765 189.515 ;
        RECT 189.620 188.965 189.970 189.175 ;
        RECT 190.140 188.965 190.585 189.165 ;
        RECT 190.755 188.965 191.230 189.165 ;
        RECT 186.890 187.975 187.220 188.435 ;
        RECT 187.730 188.145 188.480 188.435 ;
        RECT 189.705 188.625 190.770 188.795 ;
        RECT 189.705 188.145 189.875 188.625 ;
        RECT 190.045 187.975 190.375 188.455 ;
        RECT 190.600 188.395 190.770 188.625 ;
        RECT 190.950 188.565 191.230 188.965 ;
        RECT 191.500 188.965 191.830 189.165 ;
        RECT 192.000 188.965 192.365 189.165 ;
        RECT 191.500 188.565 191.785 188.965 ;
        RECT 192.595 188.795 192.765 189.345 ;
        RECT 191.965 188.625 192.765 188.795 ;
        RECT 191.965 188.395 192.135 188.625 ;
        RECT 192.935 188.555 193.105 189.685 ;
        RECT 193.295 189.435 195.885 190.525 ;
        RECT 197.010 189.725 197.260 190.525 ;
        RECT 197.430 189.895 197.760 190.355 ;
        RECT 197.930 190.065 198.145 190.525 ;
        RECT 197.430 189.725 198.600 189.895 ;
        RECT 192.920 188.475 193.105 188.555 ;
        RECT 190.600 188.145 192.135 188.395 ;
        RECT 192.305 187.975 192.635 188.455 ;
        RECT 192.850 188.145 193.105 188.475 ;
        RECT 193.295 188.745 194.505 189.265 ;
        RECT 194.675 188.915 195.885 189.435 ;
        RECT 196.520 189.555 196.800 189.715 ;
        RECT 196.520 189.385 197.855 189.555 ;
        RECT 197.685 189.215 197.855 189.385 ;
        RECT 196.520 188.965 196.870 189.205 ;
        RECT 197.040 188.965 197.515 189.205 ;
        RECT 197.685 188.965 198.060 189.215 ;
        RECT 197.685 188.795 197.855 188.965 ;
        RECT 193.295 187.975 195.885 188.745 ;
        RECT 196.520 188.625 197.855 188.795 ;
        RECT 196.520 188.415 196.790 188.625 ;
        RECT 198.230 188.435 198.600 189.725 ;
        RECT 198.815 189.435 202.325 190.525 ;
        RECT 202.495 189.435 203.705 190.525 ;
        RECT 197.010 187.975 197.340 188.435 ;
        RECT 197.850 188.145 198.600 188.435 ;
        RECT 198.815 188.745 200.465 189.265 ;
        RECT 200.635 188.915 202.325 189.435 ;
        RECT 198.815 187.975 202.325 188.745 ;
        RECT 202.495 188.725 203.015 189.265 ;
        RECT 203.185 188.895 203.705 189.435 ;
        RECT 203.875 189.360 204.165 190.525 ;
        RECT 204.335 190.090 209.680 190.525 ;
        RECT 209.855 190.090 215.200 190.525 ;
        RECT 202.495 187.975 203.705 188.725 ;
        RECT 203.875 187.975 204.165 188.700 ;
        RECT 205.920 188.520 206.260 189.350 ;
        RECT 207.740 188.840 208.090 190.090 ;
        RECT 211.440 188.520 211.780 189.350 ;
        RECT 213.260 188.840 213.610 190.090 ;
        RECT 216.295 188.920 216.575 190.355 ;
        RECT 216.745 189.750 217.455 190.525 ;
        RECT 217.625 189.580 217.955 190.355 ;
        RECT 216.805 189.365 217.955 189.580 ;
        RECT 204.335 187.975 209.680 188.520 ;
        RECT 209.855 187.975 215.200 188.520 ;
        RECT 216.295 188.145 216.635 188.920 ;
        RECT 216.805 188.795 217.090 189.365 ;
        RECT 217.275 188.965 217.745 189.195 ;
        RECT 218.150 189.165 218.365 190.280 ;
        RECT 218.545 189.805 218.875 190.525 ;
        RECT 219.055 190.090 224.400 190.525 ;
        RECT 218.655 189.165 218.885 189.505 ;
        RECT 217.915 188.985 218.365 189.165 ;
        RECT 217.915 188.965 218.245 188.985 ;
        RECT 218.555 188.965 218.885 189.165 ;
        RECT 216.805 188.605 217.515 188.795 ;
        RECT 217.215 188.465 217.515 188.605 ;
        RECT 217.705 188.605 218.885 188.795 ;
        RECT 217.705 188.525 218.035 188.605 ;
        RECT 217.215 188.455 217.530 188.465 ;
        RECT 217.215 188.445 217.540 188.455 ;
        RECT 217.215 188.440 217.550 188.445 ;
        RECT 216.805 187.975 216.975 188.435 ;
        RECT 217.215 188.430 217.555 188.440 ;
        RECT 217.215 188.425 217.560 188.430 ;
        RECT 217.215 188.415 217.565 188.425 ;
        RECT 217.215 188.410 217.570 188.415 ;
        RECT 217.215 188.145 217.575 188.410 ;
        RECT 218.205 187.975 218.375 188.435 ;
        RECT 218.545 188.145 218.885 188.605 ;
        RECT 220.640 188.520 220.980 189.350 ;
        RECT 222.460 188.840 222.810 190.090 ;
        RECT 224.575 189.435 226.245 190.525 ;
        RECT 224.575 188.745 225.325 189.265 ;
        RECT 225.495 188.915 226.245 189.435 ;
        RECT 226.415 188.920 226.695 190.355 ;
        RECT 226.865 189.750 227.575 190.525 ;
        RECT 227.745 189.580 228.075 190.355 ;
        RECT 226.925 189.365 228.075 189.580 ;
        RECT 219.055 187.975 224.400 188.520 ;
        RECT 224.575 187.975 226.245 188.745 ;
        RECT 226.415 188.145 226.755 188.920 ;
        RECT 226.925 188.795 227.210 189.365 ;
        RECT 227.395 188.965 227.865 189.195 ;
        RECT 228.270 189.165 228.485 190.280 ;
        RECT 228.665 189.805 228.995 190.525 ;
        RECT 228.775 189.165 229.005 189.505 ;
        RECT 229.635 189.360 229.925 190.525 ;
        RECT 230.185 189.595 230.355 190.355 ;
        RECT 230.535 189.765 230.865 190.525 ;
        RECT 230.185 189.425 230.850 189.595 ;
        RECT 231.035 189.450 231.305 190.355 ;
        RECT 230.680 189.280 230.850 189.425 ;
        RECT 228.035 188.985 228.485 189.165 ;
        RECT 228.035 188.965 228.365 188.985 ;
        RECT 228.675 188.965 229.005 189.165 ;
        RECT 230.115 188.875 230.445 189.245 ;
        RECT 230.680 188.950 230.965 189.280 ;
        RECT 226.925 188.605 227.635 188.795 ;
        RECT 227.335 188.465 227.635 188.605 ;
        RECT 227.825 188.605 229.005 188.795 ;
        RECT 227.825 188.525 228.155 188.605 ;
        RECT 227.335 188.455 227.650 188.465 ;
        RECT 227.335 188.445 227.660 188.455 ;
        RECT 227.335 188.440 227.670 188.445 ;
        RECT 226.925 187.975 227.095 188.435 ;
        RECT 227.335 188.430 227.675 188.440 ;
        RECT 227.335 188.425 227.680 188.430 ;
        RECT 227.335 188.415 227.685 188.425 ;
        RECT 227.335 188.410 227.690 188.415 ;
        RECT 227.335 188.145 227.695 188.410 ;
        RECT 228.325 187.975 228.495 188.435 ;
        RECT 228.665 188.145 229.005 188.605 ;
        RECT 229.635 187.975 229.925 188.700 ;
        RECT 230.680 188.695 230.850 188.950 ;
        RECT 230.185 188.525 230.850 188.695 ;
        RECT 231.135 188.650 231.305 189.450 ;
        RECT 230.185 188.145 230.355 188.525 ;
        RECT 230.535 187.975 230.865 188.355 ;
        RECT 231.045 188.145 231.305 188.650 ;
        RECT 231.475 189.450 231.745 190.355 ;
        RECT 231.915 189.765 232.245 190.525 ;
        RECT 232.425 189.595 232.595 190.355 ;
        RECT 231.475 188.650 231.645 189.450 ;
        RECT 231.930 189.425 232.595 189.595 ;
        RECT 232.855 189.450 233.125 190.355 ;
        RECT 233.295 189.765 233.625 190.525 ;
        RECT 233.805 189.595 233.975 190.355 ;
        RECT 231.930 189.280 232.100 189.425 ;
        RECT 231.815 188.950 232.100 189.280 ;
        RECT 231.930 188.695 232.100 188.950 ;
        RECT 232.335 188.875 232.665 189.245 ;
        RECT 231.475 188.145 231.735 188.650 ;
        RECT 231.930 188.525 232.595 188.695 ;
        RECT 231.915 187.975 232.245 188.355 ;
        RECT 232.425 188.145 232.595 188.525 ;
        RECT 232.855 188.650 233.025 189.450 ;
        RECT 233.310 189.425 233.975 189.595 ;
        RECT 234.235 189.435 237.745 190.525 ;
        RECT 233.310 189.280 233.480 189.425 ;
        RECT 233.195 188.950 233.480 189.280 ;
        RECT 233.310 188.695 233.480 188.950 ;
        RECT 233.715 188.875 234.045 189.245 ;
        RECT 234.235 188.745 235.885 189.265 ;
        RECT 236.055 188.915 237.745 189.435 ;
        RECT 237.915 189.435 239.125 190.525 ;
        RECT 237.915 188.895 238.435 189.435 ;
        RECT 232.855 188.145 233.115 188.650 ;
        RECT 233.310 188.525 233.975 188.695 ;
        RECT 233.295 187.975 233.625 188.355 ;
        RECT 233.805 188.145 233.975 188.525 ;
        RECT 234.235 187.975 237.745 188.745 ;
        RECT 238.605 188.725 239.125 189.265 ;
        RECT 237.915 187.975 239.125 188.725 ;
        RECT 165.150 187.805 239.210 187.975 ;
        RECT 165.235 187.055 166.445 187.805 ;
        RECT 167.165 187.255 167.335 187.635 ;
        RECT 167.515 187.425 167.845 187.805 ;
        RECT 167.165 187.085 167.830 187.255 ;
        RECT 168.025 187.130 168.285 187.635 ;
        RECT 165.235 186.515 165.755 187.055 ;
        RECT 165.925 186.345 166.445 186.885 ;
        RECT 167.095 186.535 167.425 186.905 ;
        RECT 167.660 186.830 167.830 187.085 ;
        RECT 167.660 186.500 167.945 186.830 ;
        RECT 167.660 186.355 167.830 186.500 ;
        RECT 165.235 185.255 166.445 186.345 ;
        RECT 167.165 186.185 167.830 186.355 ;
        RECT 168.115 186.330 168.285 187.130 ;
        RECT 168.545 187.255 168.715 187.635 ;
        RECT 168.895 187.425 169.225 187.805 ;
        RECT 168.545 187.085 169.210 187.255 ;
        RECT 169.405 187.130 169.665 187.635 ;
        RECT 168.475 186.535 168.805 186.905 ;
        RECT 169.040 186.830 169.210 187.085 ;
        RECT 169.040 186.500 169.325 186.830 ;
        RECT 169.040 186.355 169.210 186.500 ;
        RECT 167.165 185.425 167.335 186.185 ;
        RECT 167.515 185.255 167.845 186.015 ;
        RECT 168.015 185.425 168.285 186.330 ;
        RECT 168.545 186.185 169.210 186.355 ;
        RECT 169.495 186.330 169.665 187.130 ;
        RECT 169.925 187.255 170.095 187.635 ;
        RECT 170.310 187.425 170.640 187.805 ;
        RECT 169.925 187.085 170.640 187.255 ;
        RECT 169.835 186.535 170.190 186.905 ;
        RECT 170.470 186.895 170.640 187.085 ;
        RECT 170.810 187.060 171.065 187.635 ;
        RECT 170.470 186.565 170.725 186.895 ;
        RECT 170.470 186.355 170.640 186.565 ;
        RECT 168.545 185.425 168.715 186.185 ;
        RECT 168.895 185.255 169.225 186.015 ;
        RECT 169.395 185.425 169.665 186.330 ;
        RECT 169.925 186.185 170.640 186.355 ;
        RECT 170.895 186.330 171.065 187.060 ;
        RECT 171.240 186.965 171.500 187.805 ;
        RECT 171.735 187.325 172.015 187.805 ;
        RECT 172.185 187.155 172.445 187.545 ;
        RECT 172.620 187.325 172.875 187.805 ;
        RECT 173.045 187.155 173.340 187.545 ;
        RECT 173.520 187.325 173.795 187.805 ;
        RECT 173.965 187.305 174.265 187.635 ;
        RECT 175.360 187.405 175.695 187.805 ;
        RECT 171.690 186.985 173.340 187.155 ;
        RECT 171.690 186.475 172.095 186.985 ;
        RECT 172.265 186.645 173.405 186.815 ;
        RECT 169.925 185.425 170.095 186.185 ;
        RECT 170.310 185.255 170.640 186.015 ;
        RECT 170.810 185.425 171.065 186.330 ;
        RECT 171.240 185.255 171.500 186.405 ;
        RECT 171.690 186.305 172.445 186.475 ;
        RECT 171.730 185.255 172.015 186.125 ;
        RECT 172.185 186.055 172.445 186.305 ;
        RECT 173.235 186.395 173.405 186.645 ;
        RECT 173.575 186.565 173.925 187.135 ;
        RECT 174.095 186.395 174.265 187.305 ;
        RECT 175.865 187.235 176.070 187.635 ;
        RECT 176.280 187.325 176.555 187.805 ;
        RECT 176.765 187.305 177.025 187.635 ;
        RECT 173.235 186.225 174.265 186.395 ;
        RECT 172.185 185.885 173.305 186.055 ;
        RECT 172.185 185.425 172.445 185.885 ;
        RECT 172.620 185.255 172.875 185.715 ;
        RECT 173.045 185.425 173.305 185.885 ;
        RECT 173.475 185.255 173.785 186.055 ;
        RECT 173.955 185.425 174.265 186.225 ;
        RECT 175.385 187.065 176.070 187.235 ;
        RECT 175.385 186.035 175.725 187.065 ;
        RECT 175.895 186.395 176.145 186.895 ;
        RECT 176.325 186.565 176.685 187.145 ;
        RECT 176.855 186.395 177.025 187.305 ;
        RECT 177.350 187.155 177.680 187.620 ;
        RECT 177.850 187.335 178.020 187.805 ;
        RECT 178.190 187.155 178.520 187.635 ;
        RECT 177.350 186.985 178.520 187.155 ;
        RECT 177.195 186.605 177.840 186.815 ;
        RECT 178.010 186.605 178.580 186.815 ;
        RECT 178.750 186.435 178.920 187.635 ;
        RECT 179.460 187.235 179.630 187.440 ;
        RECT 175.895 186.225 177.025 186.395 ;
        RECT 175.385 185.860 176.050 186.035 ;
        RECT 175.360 185.255 175.695 185.680 ;
        RECT 175.865 185.455 176.050 185.860 ;
        RECT 176.255 185.255 176.585 186.035 ;
        RECT 176.755 185.455 177.025 186.225 ;
        RECT 177.410 185.255 177.740 186.355 ;
        RECT 178.215 186.025 178.920 186.435 ;
        RECT 179.090 187.065 179.630 187.235 ;
        RECT 179.910 187.065 180.080 187.805 ;
        RECT 180.345 187.065 180.705 187.440 ;
        RECT 181.425 187.255 181.595 187.635 ;
        RECT 181.775 187.425 182.105 187.805 ;
        RECT 181.425 187.085 182.090 187.255 ;
        RECT 182.285 187.130 182.545 187.635 ;
        RECT 179.090 186.365 179.260 187.065 ;
        RECT 179.430 186.565 179.760 186.895 ;
        RECT 179.930 186.565 180.280 186.895 ;
        RECT 179.090 186.195 179.715 186.365 ;
        RECT 179.930 186.025 180.195 186.565 ;
        RECT 180.450 186.410 180.705 187.065 ;
        RECT 181.355 186.535 181.685 186.905 ;
        RECT 181.920 186.830 182.090 187.085 ;
        RECT 178.215 185.855 180.195 186.025 ;
        RECT 178.215 185.425 178.540 185.855 ;
        RECT 178.710 185.255 179.040 185.675 ;
        RECT 179.785 185.255 180.195 185.685 ;
        RECT 180.365 185.425 180.705 186.410 ;
        RECT 181.920 186.500 182.205 186.830 ;
        RECT 181.920 186.355 182.090 186.500 ;
        RECT 181.425 186.185 182.090 186.355 ;
        RECT 182.375 186.330 182.545 187.130 ;
        RECT 182.805 187.255 182.975 187.635 ;
        RECT 183.155 187.425 183.485 187.805 ;
        RECT 182.805 187.085 183.470 187.255 ;
        RECT 183.665 187.130 183.925 187.635 ;
        RECT 182.735 186.535 183.065 186.905 ;
        RECT 183.300 186.830 183.470 187.085 ;
        RECT 183.300 186.500 183.585 186.830 ;
        RECT 183.300 186.355 183.470 186.500 ;
        RECT 181.425 185.425 181.595 186.185 ;
        RECT 181.775 185.255 182.105 186.015 ;
        RECT 182.275 185.425 182.545 186.330 ;
        RECT 182.805 186.185 183.470 186.355 ;
        RECT 183.755 186.330 183.925 187.130 ;
        RECT 182.805 185.425 182.975 186.185 ;
        RECT 183.155 185.255 183.485 186.015 ;
        RECT 183.655 185.425 183.925 186.330 ;
        RECT 184.095 187.130 184.355 187.635 ;
        RECT 184.535 187.425 184.865 187.805 ;
        RECT 185.045 187.255 185.215 187.635 ;
        RECT 184.095 186.330 184.265 187.130 ;
        RECT 184.550 187.085 185.215 187.255 ;
        RECT 185.565 187.255 185.735 187.635 ;
        RECT 185.915 187.425 186.245 187.805 ;
        RECT 185.565 187.085 186.230 187.255 ;
        RECT 186.425 187.130 186.685 187.635 ;
        RECT 184.550 186.830 184.720 187.085 ;
        RECT 184.435 186.500 184.720 186.830 ;
        RECT 184.955 186.535 185.285 186.905 ;
        RECT 185.495 186.535 185.825 186.905 ;
        RECT 186.060 186.830 186.230 187.085 ;
        RECT 184.550 186.355 184.720 186.500 ;
        RECT 186.060 186.500 186.345 186.830 ;
        RECT 186.060 186.355 186.230 186.500 ;
        RECT 184.095 185.425 184.365 186.330 ;
        RECT 184.550 186.185 185.215 186.355 ;
        RECT 184.535 185.255 184.865 186.015 ;
        RECT 185.045 185.425 185.215 186.185 ;
        RECT 185.565 186.185 186.230 186.355 ;
        RECT 186.515 186.330 186.685 187.130 ;
        RECT 185.565 185.425 185.735 186.185 ;
        RECT 185.915 185.255 186.245 186.015 ;
        RECT 186.415 185.425 186.685 186.330 ;
        RECT 186.855 187.130 187.115 187.635 ;
        RECT 187.295 187.425 187.625 187.805 ;
        RECT 187.805 187.255 187.975 187.635 ;
        RECT 186.855 186.330 187.025 187.130 ;
        RECT 187.310 187.085 187.975 187.255 ;
        RECT 188.235 187.130 188.495 187.635 ;
        RECT 188.675 187.425 189.005 187.805 ;
        RECT 189.185 187.255 189.355 187.635 ;
        RECT 187.310 186.830 187.480 187.085 ;
        RECT 187.195 186.500 187.480 186.830 ;
        RECT 187.715 186.535 188.045 186.905 ;
        RECT 187.310 186.355 187.480 186.500 ;
        RECT 186.855 185.425 187.125 186.330 ;
        RECT 187.310 186.185 187.975 186.355 ;
        RECT 187.295 185.255 187.625 186.015 ;
        RECT 187.805 185.425 187.975 186.185 ;
        RECT 188.235 186.330 188.405 187.130 ;
        RECT 188.690 187.085 189.355 187.255 ;
        RECT 189.615 187.130 189.875 187.635 ;
        RECT 190.055 187.425 190.385 187.805 ;
        RECT 190.565 187.255 190.735 187.635 ;
        RECT 188.690 186.830 188.860 187.085 ;
        RECT 188.575 186.500 188.860 186.830 ;
        RECT 189.095 186.535 189.425 186.905 ;
        RECT 188.690 186.355 188.860 186.500 ;
        RECT 188.235 185.425 188.505 186.330 ;
        RECT 188.690 186.185 189.355 186.355 ;
        RECT 188.675 185.255 189.005 186.015 ;
        RECT 189.185 185.425 189.355 186.185 ;
        RECT 189.615 186.330 189.785 187.130 ;
        RECT 190.070 187.085 190.735 187.255 ;
        RECT 190.070 186.830 190.240 187.085 ;
        RECT 190.995 187.080 191.285 187.805 ;
        RECT 192.005 187.255 192.175 187.635 ;
        RECT 192.355 187.425 192.685 187.805 ;
        RECT 192.005 187.085 192.670 187.255 ;
        RECT 192.865 187.130 193.125 187.635 ;
        RECT 189.955 186.500 190.240 186.830 ;
        RECT 190.475 186.535 190.805 186.905 ;
        RECT 191.935 186.535 192.265 186.905 ;
        RECT 192.500 186.830 192.670 187.085 ;
        RECT 190.070 186.355 190.240 186.500 ;
        RECT 192.500 186.500 192.785 186.830 ;
        RECT 189.615 185.425 189.885 186.330 ;
        RECT 190.070 186.185 190.735 186.355 ;
        RECT 190.055 185.255 190.385 186.015 ;
        RECT 190.565 185.425 190.735 186.185 ;
        RECT 190.995 185.255 191.285 186.420 ;
        RECT 192.500 186.355 192.670 186.500 ;
        RECT 192.005 186.185 192.670 186.355 ;
        RECT 192.955 186.330 193.125 187.130 ;
        RECT 193.845 187.155 194.015 187.635 ;
        RECT 194.185 187.325 194.515 187.805 ;
        RECT 194.740 187.385 196.275 187.635 ;
        RECT 194.740 187.155 194.910 187.385 ;
        RECT 193.845 186.985 194.910 187.155 ;
        RECT 195.090 186.815 195.370 187.215 ;
        RECT 193.760 186.605 194.110 186.815 ;
        RECT 194.280 186.615 194.725 186.815 ;
        RECT 194.895 186.615 195.370 186.815 ;
        RECT 195.640 186.815 195.925 187.215 ;
        RECT 196.105 187.155 196.275 187.385 ;
        RECT 196.445 187.325 196.775 187.805 ;
        RECT 196.990 187.305 197.245 187.635 ;
        RECT 197.060 187.225 197.245 187.305 ;
        RECT 196.105 186.985 196.905 187.155 ;
        RECT 195.640 186.615 195.970 186.815 ;
        RECT 196.140 186.615 196.505 186.815 ;
        RECT 196.735 186.435 196.905 186.985 ;
        RECT 192.005 185.425 192.175 186.185 ;
        RECT 192.355 185.255 192.685 186.015 ;
        RECT 192.855 185.425 193.125 186.330 ;
        RECT 193.845 186.265 196.905 186.435 ;
        RECT 193.845 185.425 194.015 186.265 ;
        RECT 197.075 186.095 197.245 187.225 ;
        RECT 197.985 187.155 198.155 187.635 ;
        RECT 198.325 187.325 198.655 187.805 ;
        RECT 198.880 187.385 200.415 187.635 ;
        RECT 198.880 187.155 199.050 187.385 ;
        RECT 197.985 186.985 199.050 187.155 ;
        RECT 199.230 186.815 199.510 187.215 ;
        RECT 197.900 186.605 198.250 186.815 ;
        RECT 198.420 186.615 198.865 186.815 ;
        RECT 199.035 186.615 199.510 186.815 ;
        RECT 199.780 186.815 200.065 187.215 ;
        RECT 200.245 187.155 200.415 187.385 ;
        RECT 200.585 187.325 200.915 187.805 ;
        RECT 201.130 187.305 201.385 187.635 ;
        RECT 201.175 187.295 201.385 187.305 ;
        RECT 201.200 187.225 201.385 187.295 ;
        RECT 200.245 186.985 201.045 187.155 ;
        RECT 199.780 186.615 200.110 186.815 ;
        RECT 200.280 186.615 200.645 186.815 ;
        RECT 200.875 186.435 201.045 186.985 ;
        RECT 194.185 185.595 194.515 186.095 ;
        RECT 194.685 185.855 196.320 186.095 ;
        RECT 194.685 185.765 194.915 185.855 ;
        RECT 195.025 185.595 195.355 185.635 ;
        RECT 194.185 185.425 195.355 185.595 ;
        RECT 195.545 185.255 195.900 185.675 ;
        RECT 196.070 185.425 196.320 185.855 ;
        RECT 196.490 185.255 196.820 186.015 ;
        RECT 196.990 185.425 197.245 186.095 ;
        RECT 197.985 186.265 201.045 186.435 ;
        RECT 197.985 185.425 198.155 186.265 ;
        RECT 201.215 186.095 201.385 187.225 ;
        RECT 198.325 185.595 198.655 186.095 ;
        RECT 198.825 185.855 200.460 186.095 ;
        RECT 198.825 185.765 199.055 185.855 ;
        RECT 199.165 185.595 199.495 185.635 ;
        RECT 198.325 185.425 199.495 185.595 ;
        RECT 199.685 185.255 200.040 185.675 ;
        RECT 200.210 185.425 200.460 185.855 ;
        RECT 200.630 185.255 200.960 186.015 ;
        RECT 201.130 185.425 201.385 186.095 ;
        RECT 201.575 187.130 201.835 187.635 ;
        RECT 202.015 187.425 202.345 187.805 ;
        RECT 202.525 187.255 202.695 187.635 ;
        RECT 201.575 186.330 201.745 187.130 ;
        RECT 202.030 187.085 202.695 187.255 ;
        RECT 202.030 186.830 202.200 187.085 ;
        RECT 202.955 187.035 206.465 187.805 ;
        RECT 206.635 187.055 207.845 187.805 ;
        RECT 201.915 186.500 202.200 186.830 ;
        RECT 202.435 186.535 202.765 186.905 ;
        RECT 202.955 186.515 204.605 187.035 ;
        RECT 202.030 186.355 202.200 186.500 ;
        RECT 201.575 185.425 201.845 186.330 ;
        RECT 202.030 186.185 202.695 186.355 ;
        RECT 204.775 186.345 206.465 186.865 ;
        RECT 206.635 186.515 207.155 187.055 ;
        RECT 207.325 186.345 207.845 186.885 ;
        RECT 202.015 185.255 202.345 186.015 ;
        RECT 202.525 185.425 202.695 186.185 ;
        RECT 202.955 185.255 206.465 186.345 ;
        RECT 206.635 185.255 207.845 186.345 ;
        RECT 208.015 186.860 208.355 187.635 ;
        RECT 208.525 187.345 208.695 187.805 ;
        RECT 208.935 187.370 209.295 187.635 ;
        RECT 208.935 187.365 209.290 187.370 ;
        RECT 208.935 187.355 209.285 187.365 ;
        RECT 208.935 187.350 209.280 187.355 ;
        RECT 208.935 187.340 209.275 187.350 ;
        RECT 209.925 187.345 210.095 187.805 ;
        RECT 208.935 187.335 209.270 187.340 ;
        RECT 208.935 187.325 209.260 187.335 ;
        RECT 208.935 187.315 209.250 187.325 ;
        RECT 208.935 187.175 209.235 187.315 ;
        RECT 208.525 186.985 209.235 187.175 ;
        RECT 209.425 187.175 209.755 187.255 ;
        RECT 210.265 187.175 210.605 187.635 ;
        RECT 209.425 186.985 210.605 187.175 ;
        RECT 210.775 187.130 211.035 187.635 ;
        RECT 211.215 187.425 211.545 187.805 ;
        RECT 211.725 187.255 211.895 187.635 ;
        RECT 208.015 185.425 208.295 186.860 ;
        RECT 208.525 186.415 208.810 186.985 ;
        RECT 208.995 186.585 209.465 186.815 ;
        RECT 209.635 186.795 209.965 186.815 ;
        RECT 209.635 186.615 210.085 186.795 ;
        RECT 210.275 186.615 210.605 186.815 ;
        RECT 208.525 186.200 209.675 186.415 ;
        RECT 208.465 185.255 209.175 186.030 ;
        RECT 209.345 185.425 209.675 186.200 ;
        RECT 209.870 185.500 210.085 186.615 ;
        RECT 210.375 186.275 210.605 186.615 ;
        RECT 210.775 186.330 210.945 187.130 ;
        RECT 211.230 187.085 211.895 187.255 ;
        RECT 212.155 187.130 212.415 187.635 ;
        RECT 212.595 187.425 212.925 187.805 ;
        RECT 213.105 187.255 213.275 187.635 ;
        RECT 211.230 186.830 211.400 187.085 ;
        RECT 211.115 186.500 211.400 186.830 ;
        RECT 211.635 186.535 211.965 186.905 ;
        RECT 211.230 186.355 211.400 186.500 ;
        RECT 210.265 185.255 210.595 185.975 ;
        RECT 210.775 185.425 211.045 186.330 ;
        RECT 211.230 186.185 211.895 186.355 ;
        RECT 211.215 185.255 211.545 186.015 ;
        RECT 211.725 185.425 211.895 186.185 ;
        RECT 212.155 186.330 212.325 187.130 ;
        RECT 212.610 187.085 213.275 187.255 ;
        RECT 213.625 187.255 213.795 187.635 ;
        RECT 213.975 187.425 214.305 187.805 ;
        RECT 213.625 187.085 214.290 187.255 ;
        RECT 214.485 187.130 214.745 187.635 ;
        RECT 212.610 186.830 212.780 187.085 ;
        RECT 212.495 186.500 212.780 186.830 ;
        RECT 213.015 186.535 213.345 186.905 ;
        RECT 213.555 186.535 213.885 186.905 ;
        RECT 214.120 186.830 214.290 187.085 ;
        RECT 212.610 186.355 212.780 186.500 ;
        RECT 214.120 186.500 214.405 186.830 ;
        RECT 214.120 186.355 214.290 186.500 ;
        RECT 212.155 185.425 212.425 186.330 ;
        RECT 212.610 186.185 213.275 186.355 ;
        RECT 212.595 185.255 212.925 186.015 ;
        RECT 213.105 185.425 213.275 186.185 ;
        RECT 213.625 186.185 214.290 186.355 ;
        RECT 214.575 186.330 214.745 187.130 ;
        RECT 215.005 187.255 215.175 187.635 ;
        RECT 215.355 187.425 215.685 187.805 ;
        RECT 215.005 187.085 215.670 187.255 ;
        RECT 215.865 187.130 216.125 187.635 ;
        RECT 214.935 186.535 215.265 186.905 ;
        RECT 215.500 186.830 215.670 187.085 ;
        RECT 215.500 186.500 215.785 186.830 ;
        RECT 215.500 186.355 215.670 186.500 ;
        RECT 213.625 185.425 213.795 186.185 ;
        RECT 213.975 185.255 214.305 186.015 ;
        RECT 214.475 185.425 214.745 186.330 ;
        RECT 215.005 186.185 215.670 186.355 ;
        RECT 215.955 186.330 216.125 187.130 ;
        RECT 216.755 187.080 217.045 187.805 ;
        RECT 217.305 187.255 217.475 187.635 ;
        RECT 217.655 187.425 217.985 187.805 ;
        RECT 217.305 187.085 217.970 187.255 ;
        RECT 218.165 187.130 218.425 187.635 ;
        RECT 217.235 186.535 217.565 186.905 ;
        RECT 217.800 186.830 217.970 187.085 ;
        RECT 217.800 186.500 218.085 186.830 ;
        RECT 215.005 185.425 215.175 186.185 ;
        RECT 215.355 185.255 215.685 186.015 ;
        RECT 215.855 185.425 216.125 186.330 ;
        RECT 216.755 185.255 217.045 186.420 ;
        RECT 217.800 186.355 217.970 186.500 ;
        RECT 217.305 186.185 217.970 186.355 ;
        RECT 218.255 186.330 218.425 187.130 ;
        RECT 218.685 187.255 218.855 187.635 ;
        RECT 219.035 187.425 219.365 187.805 ;
        RECT 218.685 187.085 219.350 187.255 ;
        RECT 219.545 187.130 219.805 187.635 ;
        RECT 218.615 186.535 218.945 186.905 ;
        RECT 219.180 186.830 219.350 187.085 ;
        RECT 219.180 186.500 219.465 186.830 ;
        RECT 219.180 186.355 219.350 186.500 ;
        RECT 217.305 185.425 217.475 186.185 ;
        RECT 217.655 185.255 217.985 186.015 ;
        RECT 218.155 185.425 218.425 186.330 ;
        RECT 218.685 186.185 219.350 186.355 ;
        RECT 219.635 186.330 219.805 187.130 ;
        RECT 218.685 185.425 218.855 186.185 ;
        RECT 219.035 185.255 219.365 186.015 ;
        RECT 219.535 185.425 219.805 186.330 ;
        RECT 219.975 187.130 220.235 187.635 ;
        RECT 220.415 187.425 220.745 187.805 ;
        RECT 220.925 187.255 221.095 187.635 ;
        RECT 219.975 186.330 220.145 187.130 ;
        RECT 220.430 187.085 221.095 187.255 ;
        RECT 221.445 187.255 221.615 187.635 ;
        RECT 221.795 187.425 222.125 187.805 ;
        RECT 221.445 187.085 222.110 187.255 ;
        RECT 222.305 187.130 222.565 187.635 ;
        RECT 220.430 186.830 220.600 187.085 ;
        RECT 220.315 186.500 220.600 186.830 ;
        RECT 220.835 186.535 221.165 186.905 ;
        RECT 221.375 186.535 221.705 186.905 ;
        RECT 221.940 186.830 222.110 187.085 ;
        RECT 220.430 186.355 220.600 186.500 ;
        RECT 221.940 186.500 222.225 186.830 ;
        RECT 221.940 186.355 222.110 186.500 ;
        RECT 219.975 185.425 220.245 186.330 ;
        RECT 220.430 186.185 221.095 186.355 ;
        RECT 220.415 185.255 220.745 186.015 ;
        RECT 220.925 185.425 221.095 186.185 ;
        RECT 221.445 186.185 222.110 186.355 ;
        RECT 222.395 186.330 222.565 187.130 ;
        RECT 222.825 187.255 222.995 187.630 ;
        RECT 223.165 187.425 223.495 187.805 ;
        RECT 223.665 187.465 224.740 187.635 ;
        RECT 223.665 187.255 223.835 187.465 ;
        RECT 222.825 187.085 223.835 187.255 ;
        RECT 224.060 187.125 224.400 187.295 ;
        RECT 224.570 187.130 224.740 187.465 ;
        RECT 224.060 186.955 224.350 187.125 ;
        RECT 222.800 186.445 223.145 186.895 ;
        RECT 221.445 185.425 221.615 186.185 ;
        RECT 221.795 185.255 222.125 186.015 ;
        RECT 222.295 185.425 222.565 186.330 ;
        RECT 222.795 186.275 223.145 186.445 ;
        RECT 223.455 186.275 223.890 186.895 ;
        RECT 224.060 186.435 224.230 186.955 ;
        RECT 224.910 186.785 225.270 187.460 ;
        RECT 225.450 187.085 225.740 187.805 ;
        RECT 226.030 187.465 227.630 187.635 ;
        RECT 226.030 187.095 226.200 187.465 ;
        RECT 227.275 187.425 227.630 187.465 ;
        RECT 227.800 187.345 227.970 187.805 ;
        RECT 226.370 187.045 226.700 187.295 ;
        RECT 226.385 186.970 226.700 187.045 ;
        RECT 226.870 187.175 227.040 187.295 ;
        RECT 228.145 187.175 228.390 187.595 ;
        RECT 228.660 187.425 228.990 187.805 ;
        RECT 229.160 187.235 229.335 187.565 ;
        RECT 229.680 187.475 229.850 187.635 ;
        RECT 229.680 187.305 230.210 187.475 ;
        RECT 230.380 187.465 231.375 187.635 ;
        RECT 230.380 187.305 230.550 187.465 ;
        RECT 226.870 187.005 228.390 187.175 ;
        RECT 224.730 186.605 225.270 186.785 ;
        RECT 224.910 186.495 225.270 186.605 ;
        RECT 224.060 186.265 224.695 186.435 ;
        RECT 224.910 186.265 225.715 186.495 ;
        RECT 222.825 185.925 224.355 186.095 ;
        RECT 222.825 185.425 222.995 185.925 ;
        RECT 224.185 185.765 224.355 185.925 ;
        RECT 224.525 185.935 224.695 186.265 ;
        RECT 224.525 185.765 224.855 185.935 ;
        RECT 223.165 185.255 223.495 185.635 ;
        RECT 223.665 185.595 223.835 185.755 ;
        RECT 225.025 185.595 225.195 186.095 ;
        RECT 223.665 185.425 225.195 185.595 ;
        RECT 225.365 185.425 225.715 186.265 ;
        RECT 225.915 185.895 226.215 186.895 ;
        RECT 226.385 186.445 226.555 186.970 ;
        RECT 226.870 186.965 227.040 187.005 ;
        RECT 226.725 186.785 227.055 186.795 ;
        RECT 226.725 186.625 227.110 186.785 ;
        RECT 226.940 186.615 227.110 186.625 ;
        RECT 227.450 186.445 227.695 186.835 ;
        RECT 226.385 186.275 227.145 186.445 ;
        RECT 227.395 186.275 227.695 186.445 ;
        RECT 225.885 185.255 226.215 185.635 ;
        RECT 226.475 185.595 226.645 186.105 ;
        RECT 226.815 185.765 227.145 186.275 ;
        RECT 227.450 186.215 227.695 186.275 ;
        RECT 227.900 186.215 228.230 186.835 ;
        RECT 228.705 186.215 228.995 186.895 ;
        RECT 229.165 186.785 229.335 187.235 ;
        RECT 229.630 186.955 229.870 187.125 ;
        RECT 229.165 186.615 229.455 186.785 ;
        RECT 227.315 185.805 228.380 185.975 ;
        RECT 227.315 185.595 227.485 185.805 ;
        RECT 226.475 185.425 227.485 185.595 ;
        RECT 227.710 185.255 228.040 185.635 ;
        RECT 228.210 185.425 228.380 185.805 ;
        RECT 229.165 185.755 229.335 186.615 ;
        RECT 228.630 185.255 228.980 185.635 ;
        RECT 229.150 185.425 229.335 185.755 ;
        RECT 229.630 185.755 229.800 186.955 ;
        RECT 230.040 186.135 230.210 187.305 ;
        RECT 230.860 187.125 231.035 187.295 ;
        RECT 230.620 186.965 231.035 187.125 ;
        RECT 231.205 187.175 231.375 187.465 ;
        RECT 231.545 187.345 231.715 187.805 ;
        RECT 231.205 187.005 231.775 187.175 ;
        RECT 230.620 186.955 231.030 186.965 ;
        RECT 230.840 186.615 231.295 186.785 ;
        RECT 231.605 186.225 231.775 187.005 ;
        RECT 230.040 185.905 230.825 186.135 ;
        RECT 230.495 185.765 230.825 185.905 ;
        RECT 231.125 186.055 231.775 186.225 ;
        RECT 229.630 185.425 229.840 185.755 ;
        RECT 230.010 185.595 230.340 185.635 ;
        RECT 231.125 185.595 231.295 186.055 ;
        RECT 230.010 185.425 231.295 185.595 ;
        RECT 231.465 185.255 231.795 185.635 ;
        RECT 231.965 185.425 232.225 187.635 ;
        RECT 232.395 187.175 232.735 187.635 ;
        RECT 232.905 187.345 233.075 187.805 ;
        RECT 233.705 187.370 234.065 187.635 ;
        RECT 233.710 187.365 234.065 187.370 ;
        RECT 233.715 187.355 234.065 187.365 ;
        RECT 233.720 187.350 234.065 187.355 ;
        RECT 233.725 187.340 234.065 187.350 ;
        RECT 234.305 187.345 234.475 187.805 ;
        RECT 233.730 187.335 234.065 187.340 ;
        RECT 233.740 187.325 234.065 187.335 ;
        RECT 233.750 187.315 234.065 187.325 ;
        RECT 233.245 187.175 233.575 187.255 ;
        RECT 232.395 186.985 233.575 187.175 ;
        RECT 233.765 187.175 234.065 187.315 ;
        RECT 233.765 186.985 234.475 187.175 ;
        RECT 232.395 186.615 232.725 186.815 ;
        RECT 233.035 186.795 233.365 186.815 ;
        RECT 232.915 186.615 233.365 186.795 ;
        RECT 232.395 186.275 232.625 186.615 ;
        RECT 232.405 185.255 232.735 185.975 ;
        RECT 232.915 185.500 233.130 186.615 ;
        RECT 233.535 186.585 234.005 186.815 ;
        RECT 234.190 186.415 234.475 186.985 ;
        RECT 234.645 186.860 234.985 187.635 ;
        RECT 233.325 186.200 234.475 186.415 ;
        RECT 233.325 185.425 233.655 186.200 ;
        RECT 233.825 185.255 234.535 186.030 ;
        RECT 234.705 185.425 234.985 186.860 ;
        RECT 235.155 187.130 235.415 187.635 ;
        RECT 235.595 187.425 235.925 187.805 ;
        RECT 236.105 187.255 236.275 187.635 ;
        RECT 235.155 186.330 235.325 187.130 ;
        RECT 235.610 187.085 236.275 187.255 ;
        RECT 235.610 186.830 235.780 187.085 ;
        RECT 236.535 187.055 237.745 187.805 ;
        RECT 237.915 187.055 239.125 187.805 ;
        RECT 235.495 186.500 235.780 186.830 ;
        RECT 236.015 186.535 236.345 186.905 ;
        RECT 236.535 186.515 237.055 187.055 ;
        RECT 235.610 186.355 235.780 186.500 ;
        RECT 235.155 185.425 235.425 186.330 ;
        RECT 235.610 186.185 236.275 186.355 ;
        RECT 237.225 186.345 237.745 186.885 ;
        RECT 235.595 185.255 235.925 186.015 ;
        RECT 236.105 185.425 236.275 186.185 ;
        RECT 236.535 185.255 237.745 186.345 ;
        RECT 237.915 186.345 238.435 186.885 ;
        RECT 238.605 186.515 239.125 187.055 ;
        RECT 237.915 185.255 239.125 186.345 ;
        RECT 165.150 185.085 239.210 185.255 ;
        RECT 108.630 184.880 153.130 185.050 ;
        RECT 165.235 183.995 166.445 185.085 ;
        RECT 165.235 183.285 165.755 183.825 ;
        RECT 165.925 183.455 166.445 183.995 ;
        RECT 166.705 184.155 166.875 184.915 ;
        RECT 167.055 184.325 167.385 185.085 ;
        RECT 166.705 183.985 167.370 184.155 ;
        RECT 167.555 184.010 167.825 184.915 ;
        RECT 167.200 183.840 167.370 183.985 ;
        RECT 166.635 183.435 166.965 183.805 ;
        RECT 167.200 183.510 167.485 183.840 ;
        RECT 165.235 182.535 166.445 183.285 ;
        RECT 167.200 183.255 167.370 183.510 ;
        RECT 166.705 183.085 167.370 183.255 ;
        RECT 167.655 183.210 167.825 184.010 ;
        RECT 168.000 183.935 168.260 185.085 ;
        RECT 168.435 184.010 168.690 184.915 ;
        RECT 168.860 184.325 169.190 185.085 ;
        RECT 169.405 184.155 169.575 184.915 ;
        RECT 166.705 182.705 166.875 183.085 ;
        RECT 167.055 182.535 167.385 182.915 ;
        RECT 167.565 182.705 167.825 183.210 ;
        RECT 168.000 182.535 168.260 183.375 ;
        RECT 168.435 183.280 168.605 184.010 ;
        RECT 168.860 183.985 169.575 184.155 ;
        RECT 169.855 184.245 170.110 184.915 ;
        RECT 170.280 184.325 170.610 185.085 ;
        RECT 170.780 184.485 171.030 184.915 ;
        RECT 171.200 184.665 171.555 185.085 ;
        RECT 171.745 184.745 172.915 184.915 ;
        RECT 171.745 184.705 172.075 184.745 ;
        RECT 172.185 184.485 172.415 184.575 ;
        RECT 170.780 184.245 172.415 184.485 ;
        RECT 172.585 184.245 172.915 184.745 ;
        RECT 168.860 183.775 169.030 183.985 ;
        RECT 168.775 183.445 169.030 183.775 ;
        RECT 168.435 182.705 168.690 183.280 ;
        RECT 168.860 183.255 169.030 183.445 ;
        RECT 169.310 183.435 169.665 183.805 ;
        RECT 168.860 183.085 169.575 183.255 ;
        RECT 168.860 182.535 169.190 182.915 ;
        RECT 169.405 182.705 169.575 183.085 ;
        RECT 169.855 183.115 170.025 184.245 ;
        RECT 173.085 184.075 173.255 184.915 ;
        RECT 170.195 183.905 173.255 184.075 ;
        RECT 174.525 184.075 174.695 184.915 ;
        RECT 174.865 184.745 176.035 184.915 ;
        RECT 174.865 184.245 175.195 184.745 ;
        RECT 175.705 184.705 176.035 184.745 ;
        RECT 176.225 184.665 176.580 185.085 ;
        RECT 175.365 184.485 175.595 184.575 ;
        RECT 176.750 184.485 177.000 184.915 ;
        RECT 175.365 184.245 177.000 184.485 ;
        RECT 177.170 184.325 177.500 185.085 ;
        RECT 177.670 184.245 177.925 184.915 ;
        RECT 174.525 183.905 177.585 184.075 ;
        RECT 170.195 183.355 170.365 183.905 ;
        RECT 170.585 183.555 170.960 183.725 ;
        RECT 170.595 183.525 170.960 183.555 ;
        RECT 171.130 183.525 171.460 183.725 ;
        RECT 170.195 183.185 170.995 183.355 ;
        RECT 169.855 183.035 170.040 183.115 ;
        RECT 169.855 182.705 170.110 183.035 ;
        RECT 170.325 182.535 170.655 183.015 ;
        RECT 170.825 182.955 170.995 183.185 ;
        RECT 171.175 183.125 171.460 183.525 ;
        RECT 171.730 183.525 172.205 183.725 ;
        RECT 172.375 183.525 172.820 183.725 ;
        RECT 172.990 183.525 173.340 183.735 ;
        RECT 174.440 183.525 174.790 183.735 ;
        RECT 174.960 183.525 175.405 183.725 ;
        RECT 175.575 183.525 176.050 183.725 ;
        RECT 171.730 183.125 172.010 183.525 ;
        RECT 172.190 183.185 173.255 183.355 ;
        RECT 172.190 182.955 172.360 183.185 ;
        RECT 170.825 182.705 172.360 182.955 ;
        RECT 172.585 182.535 172.915 183.015 ;
        RECT 173.085 182.705 173.255 183.185 ;
        RECT 174.525 183.185 175.590 183.355 ;
        RECT 174.525 182.705 174.695 183.185 ;
        RECT 174.865 182.535 175.195 183.015 ;
        RECT 175.420 182.955 175.590 183.185 ;
        RECT 175.770 183.125 176.050 183.525 ;
        RECT 176.320 183.525 176.650 183.725 ;
        RECT 176.820 183.555 177.195 183.725 ;
        RECT 176.820 183.525 177.185 183.555 ;
        RECT 176.320 183.125 176.605 183.525 ;
        RECT 177.415 183.355 177.585 183.905 ;
        RECT 176.785 183.185 177.585 183.355 ;
        RECT 176.785 182.955 176.955 183.185 ;
        RECT 177.755 183.115 177.925 184.245 ;
        RECT 178.115 183.920 178.405 185.085 ;
        RECT 178.790 183.985 179.120 185.085 ;
        RECT 179.595 184.485 179.920 184.915 ;
        RECT 180.090 184.665 180.420 185.085 ;
        RECT 181.165 184.655 181.575 185.085 ;
        RECT 179.595 184.315 181.575 184.485 ;
        RECT 179.595 183.905 180.300 184.315 ;
        RECT 178.575 183.525 179.220 183.735 ;
        RECT 179.390 183.525 179.960 183.735 ;
        RECT 177.740 183.035 177.925 183.115 ;
        RECT 175.420 182.705 176.955 182.955 ;
        RECT 177.125 182.535 177.455 183.015 ;
        RECT 177.670 182.705 177.925 183.035 ;
        RECT 178.115 182.535 178.405 183.260 ;
        RECT 178.730 183.185 179.900 183.355 ;
        RECT 178.730 182.720 179.060 183.185 ;
        RECT 179.230 182.535 179.400 183.005 ;
        RECT 179.570 182.705 179.900 183.185 ;
        RECT 180.130 182.705 180.300 183.905 ;
        RECT 180.470 183.975 181.095 184.145 ;
        RECT 180.470 183.275 180.640 183.975 ;
        RECT 181.310 183.775 181.575 184.315 ;
        RECT 181.745 183.930 182.085 184.915 ;
        RECT 182.805 184.155 182.975 184.915 ;
        RECT 183.155 184.325 183.485 185.085 ;
        RECT 182.805 183.985 183.470 184.155 ;
        RECT 183.655 184.010 183.925 184.915 ;
        RECT 184.590 184.285 184.840 185.085 ;
        RECT 185.010 184.455 185.340 184.915 ;
        RECT 185.510 184.625 185.725 185.085 ;
        RECT 185.010 184.285 186.180 184.455 ;
        RECT 186.890 184.285 187.140 185.085 ;
        RECT 187.310 184.455 187.640 184.915 ;
        RECT 187.810 184.625 188.025 185.085 ;
        RECT 187.310 184.285 188.480 184.455 ;
        RECT 180.810 183.445 181.140 183.775 ;
        RECT 181.310 183.445 181.660 183.775 ;
        RECT 181.830 183.275 182.085 183.930 ;
        RECT 183.300 183.840 183.470 183.985 ;
        RECT 182.735 183.435 183.065 183.805 ;
        RECT 183.300 183.510 183.585 183.840 ;
        RECT 180.470 183.105 181.010 183.275 ;
        RECT 180.840 182.900 181.010 183.105 ;
        RECT 181.290 182.535 181.460 183.275 ;
        RECT 181.725 182.900 182.085 183.275 ;
        RECT 183.300 183.255 183.470 183.510 ;
        RECT 182.805 183.085 183.470 183.255 ;
        RECT 183.755 183.210 183.925 184.010 ;
        RECT 184.100 184.115 184.380 184.275 ;
        RECT 184.100 183.945 185.435 184.115 ;
        RECT 185.265 183.775 185.435 183.945 ;
        RECT 184.100 183.525 184.450 183.765 ;
        RECT 184.620 183.525 185.095 183.765 ;
        RECT 185.265 183.525 185.640 183.775 ;
        RECT 185.265 183.355 185.435 183.525 ;
        RECT 182.805 182.705 182.975 183.085 ;
        RECT 183.155 182.535 183.485 182.915 ;
        RECT 183.665 182.705 183.925 183.210 ;
        RECT 184.100 183.185 185.435 183.355 ;
        RECT 184.100 182.975 184.370 183.185 ;
        RECT 185.810 182.995 186.180 184.285 ;
        RECT 186.400 184.115 186.680 184.275 ;
        RECT 186.400 183.945 187.735 184.115 ;
        RECT 187.565 183.775 187.735 183.945 ;
        RECT 186.400 183.525 186.750 183.765 ;
        RECT 186.920 183.525 187.395 183.765 ;
        RECT 187.565 183.525 187.940 183.775 ;
        RECT 187.565 183.355 187.735 183.525 ;
        RECT 184.590 182.535 184.920 182.995 ;
        RECT 185.430 182.705 186.180 182.995 ;
        RECT 186.400 183.185 187.735 183.355 ;
        RECT 186.400 182.975 186.670 183.185 ;
        RECT 188.110 182.995 188.480 184.285 ;
        RECT 188.785 184.075 188.955 184.915 ;
        RECT 189.125 184.745 190.295 184.915 ;
        RECT 189.125 184.245 189.455 184.745 ;
        RECT 189.965 184.705 190.295 184.745 ;
        RECT 190.485 184.665 190.840 185.085 ;
        RECT 189.625 184.485 189.855 184.575 ;
        RECT 191.010 184.485 191.260 184.915 ;
        RECT 189.625 184.245 191.260 184.485 ;
        RECT 191.430 184.325 191.760 185.085 ;
        RECT 191.930 184.245 192.185 184.915 ;
        RECT 188.785 183.905 191.845 184.075 ;
        RECT 188.700 183.525 189.050 183.735 ;
        RECT 189.220 183.525 189.665 183.725 ;
        RECT 189.835 183.525 190.310 183.725 ;
        RECT 186.890 182.535 187.220 182.995 ;
        RECT 187.730 182.705 188.480 182.995 ;
        RECT 188.785 183.185 189.850 183.355 ;
        RECT 188.785 182.705 188.955 183.185 ;
        RECT 189.125 182.535 189.455 183.015 ;
        RECT 189.680 182.955 189.850 183.185 ;
        RECT 190.030 183.125 190.310 183.525 ;
        RECT 190.580 183.525 190.910 183.725 ;
        RECT 191.080 183.525 191.445 183.725 ;
        RECT 190.580 183.125 190.865 183.525 ;
        RECT 191.675 183.355 191.845 183.905 ;
        RECT 191.045 183.185 191.845 183.355 ;
        RECT 191.045 182.955 191.215 183.185 ;
        RECT 192.015 183.115 192.185 184.245 ;
        RECT 192.000 183.045 192.185 183.115 ;
        RECT 191.975 183.035 192.185 183.045 ;
        RECT 189.680 182.705 191.215 182.955 ;
        RECT 191.385 182.535 191.715 183.015 ;
        RECT 191.930 182.705 192.185 183.035 ;
        RECT 192.380 183.945 192.715 184.915 ;
        RECT 192.885 183.945 193.055 185.085 ;
        RECT 193.225 184.745 195.255 184.915 ;
        RECT 192.380 183.275 192.550 183.945 ;
        RECT 193.225 183.775 193.395 184.745 ;
        RECT 192.720 183.445 192.975 183.775 ;
        RECT 193.200 183.445 193.395 183.775 ;
        RECT 193.565 184.405 194.690 184.575 ;
        RECT 192.805 183.275 192.975 183.445 ;
        RECT 193.565 183.275 193.735 184.405 ;
        RECT 192.380 182.705 192.635 183.275 ;
        RECT 192.805 183.105 193.735 183.275 ;
        RECT 193.905 184.065 194.915 184.235 ;
        RECT 193.905 183.265 194.075 184.065 ;
        RECT 193.560 183.070 193.735 183.105 ;
        RECT 192.805 182.535 193.135 182.935 ;
        RECT 193.560 182.705 194.090 183.070 ;
        RECT 194.280 183.045 194.555 183.865 ;
        RECT 194.275 182.875 194.555 183.045 ;
        RECT 194.280 182.705 194.555 182.875 ;
        RECT 194.725 182.705 194.915 184.065 ;
        RECT 195.085 184.080 195.255 184.745 ;
        RECT 195.425 184.325 195.595 185.085 ;
        RECT 195.830 184.325 196.345 184.735 ;
        RECT 195.085 183.890 195.835 184.080 ;
        RECT 196.005 183.515 196.345 184.325 ;
        RECT 197.065 184.075 197.235 184.915 ;
        RECT 197.405 184.745 198.575 184.915 ;
        RECT 197.405 184.245 197.735 184.745 ;
        RECT 198.245 184.705 198.575 184.745 ;
        RECT 198.765 184.665 199.120 185.085 ;
        RECT 197.905 184.485 198.135 184.575 ;
        RECT 199.290 184.485 199.540 184.915 ;
        RECT 197.905 184.245 199.540 184.485 ;
        RECT 199.710 184.325 200.040 185.085 ;
        RECT 200.210 184.245 200.465 184.915 ;
        RECT 200.255 184.235 200.465 184.245 ;
        RECT 197.065 183.905 200.125 184.075 ;
        RECT 196.980 183.525 197.330 183.735 ;
        RECT 197.500 183.525 197.945 183.725 ;
        RECT 198.115 183.525 198.590 183.725 ;
        RECT 195.115 183.345 196.345 183.515 ;
        RECT 195.095 182.535 195.605 183.070 ;
        RECT 195.825 182.740 196.070 183.345 ;
        RECT 197.065 183.185 198.130 183.355 ;
        RECT 197.065 182.705 197.235 183.185 ;
        RECT 197.405 182.535 197.735 183.015 ;
        RECT 197.960 182.955 198.130 183.185 ;
        RECT 198.310 183.125 198.590 183.525 ;
        RECT 198.860 183.525 199.190 183.725 ;
        RECT 199.360 183.525 199.725 183.725 ;
        RECT 198.860 183.125 199.145 183.525 ;
        RECT 199.955 183.355 200.125 183.905 ;
        RECT 199.325 183.185 200.125 183.355 ;
        RECT 199.325 182.955 199.495 183.185 ;
        RECT 200.295 183.115 200.465 184.235 ;
        RECT 200.280 183.035 200.465 183.115 ;
        RECT 197.960 182.705 199.495 182.955 ;
        RECT 199.665 182.535 199.995 183.015 ;
        RECT 200.210 182.705 200.465 183.035 ;
        RECT 201.115 184.010 201.385 184.915 ;
        RECT 201.555 184.325 201.885 185.085 ;
        RECT 202.065 184.155 202.235 184.915 ;
        RECT 201.115 183.210 201.285 184.010 ;
        RECT 201.570 183.985 202.235 184.155 ;
        RECT 202.495 184.010 202.765 184.915 ;
        RECT 202.935 184.325 203.265 185.085 ;
        RECT 203.445 184.155 203.615 184.915 ;
        RECT 201.570 183.840 201.740 183.985 ;
        RECT 201.455 183.510 201.740 183.840 ;
        RECT 201.570 183.255 201.740 183.510 ;
        RECT 201.975 183.435 202.305 183.805 ;
        RECT 201.115 182.705 201.375 183.210 ;
        RECT 201.570 183.085 202.235 183.255 ;
        RECT 201.555 182.535 201.885 182.915 ;
        RECT 202.065 182.705 202.235 183.085 ;
        RECT 202.495 183.210 202.665 184.010 ;
        RECT 202.950 183.985 203.615 184.155 ;
        RECT 202.950 183.840 203.120 183.985 ;
        RECT 203.875 183.920 204.165 185.085 ;
        RECT 204.335 183.995 206.005 185.085 ;
        RECT 202.835 183.510 203.120 183.840 ;
        RECT 202.950 183.255 203.120 183.510 ;
        RECT 203.355 183.435 203.685 183.805 ;
        RECT 204.335 183.305 205.085 183.825 ;
        RECT 205.255 183.475 206.005 183.995 ;
        RECT 206.725 184.155 206.895 184.915 ;
        RECT 207.075 184.325 207.405 185.085 ;
        RECT 206.725 183.985 207.390 184.155 ;
        RECT 207.575 184.010 207.845 184.915 ;
        RECT 208.105 184.415 208.275 184.915 ;
        RECT 208.445 184.705 208.775 185.085 ;
        RECT 208.945 184.745 210.475 184.915 ;
        RECT 208.945 184.585 209.115 184.745 ;
        RECT 209.465 184.415 209.635 184.575 ;
        RECT 208.105 184.245 209.635 184.415 ;
        RECT 209.805 184.405 210.135 184.575 ;
        RECT 209.805 184.075 209.975 184.405 ;
        RECT 210.305 184.245 210.475 184.745 ;
        RECT 210.645 184.075 210.995 184.915 ;
        RECT 211.165 184.705 211.495 185.085 ;
        RECT 211.755 184.745 212.765 184.915 ;
        RECT 207.220 183.840 207.390 183.985 ;
        RECT 206.655 183.435 206.985 183.805 ;
        RECT 207.220 183.510 207.505 183.840 ;
        RECT 202.495 182.705 202.755 183.210 ;
        RECT 202.950 183.085 203.615 183.255 ;
        RECT 202.935 182.535 203.265 182.915 ;
        RECT 203.445 182.705 203.615 183.085 ;
        RECT 203.875 182.535 204.165 183.260 ;
        RECT 204.335 182.535 206.005 183.305 ;
        RECT 207.220 183.255 207.390 183.510 ;
        RECT 206.725 183.085 207.390 183.255 ;
        RECT 207.675 183.210 207.845 184.010 ;
        RECT 208.075 183.895 208.425 184.065 ;
        RECT 208.080 183.445 208.425 183.895 ;
        RECT 208.735 183.445 209.170 184.065 ;
        RECT 209.340 183.905 209.975 184.075 ;
        RECT 209.340 183.385 209.510 183.905 ;
        RECT 210.190 183.845 210.995 184.075 ;
        RECT 210.190 183.735 210.550 183.845 ;
        RECT 210.010 183.555 210.550 183.735 ;
        RECT 206.725 182.705 206.895 183.085 ;
        RECT 207.075 182.535 207.405 182.915 ;
        RECT 207.585 182.705 207.845 183.210 ;
        RECT 208.105 183.085 209.115 183.255 ;
        RECT 208.105 182.710 208.275 183.085 ;
        RECT 208.445 182.535 208.775 182.915 ;
        RECT 208.945 182.875 209.115 183.085 ;
        RECT 209.340 183.215 209.630 183.385 ;
        RECT 209.340 183.045 209.680 183.215 ;
        RECT 209.850 182.875 210.020 183.210 ;
        RECT 210.190 182.880 210.550 183.555 ;
        RECT 211.195 183.445 211.495 184.445 ;
        RECT 211.755 184.235 211.925 184.745 ;
        RECT 212.095 184.065 212.425 184.575 ;
        RECT 212.595 184.535 212.765 184.745 ;
        RECT 212.990 184.705 213.320 185.085 ;
        RECT 213.490 184.535 213.660 184.915 ;
        RECT 213.910 184.705 214.260 185.085 ;
        RECT 214.430 184.585 214.615 184.915 ;
        RECT 212.595 184.365 213.660 184.535 ;
        RECT 212.730 184.065 212.975 184.125 ;
        RECT 211.665 183.895 212.425 184.065 ;
        RECT 212.675 183.895 212.975 184.065 ;
        RECT 211.665 183.370 211.835 183.895 ;
        RECT 212.220 183.715 212.390 183.725 ;
        RECT 212.005 183.555 212.390 183.715 ;
        RECT 212.005 183.545 212.335 183.555 ;
        RECT 212.730 183.505 212.975 183.895 ;
        RECT 213.180 183.505 213.510 184.125 ;
        RECT 213.985 183.445 214.275 184.125 ;
        RECT 214.445 183.725 214.615 184.585 ;
        RECT 214.910 184.585 215.120 184.915 ;
        RECT 215.290 184.745 216.575 184.915 ;
        RECT 215.290 184.705 215.620 184.745 ;
        RECT 214.445 183.555 214.735 183.725 ;
        RECT 211.665 183.295 211.980 183.370 ;
        RECT 208.945 182.705 210.020 182.875 ;
        RECT 210.730 182.535 211.020 183.255 ;
        RECT 211.310 182.875 211.480 183.245 ;
        RECT 211.650 183.045 211.980 183.295 ;
        RECT 212.150 183.335 212.320 183.375 ;
        RECT 212.150 183.165 213.670 183.335 ;
        RECT 212.150 183.045 212.320 183.165 ;
        RECT 212.555 182.875 212.910 182.915 ;
        RECT 211.310 182.705 212.910 182.875 ;
        RECT 213.080 182.535 213.250 182.995 ;
        RECT 213.425 182.745 213.670 183.165 ;
        RECT 214.445 183.105 214.615 183.555 ;
        RECT 214.910 183.385 215.080 184.585 ;
        RECT 215.775 184.435 216.105 184.575 ;
        RECT 215.320 184.205 216.105 184.435 ;
        RECT 216.405 184.285 216.575 184.745 ;
        RECT 216.745 184.705 217.075 185.085 ;
        RECT 214.910 183.215 215.150 183.385 ;
        RECT 213.940 182.535 214.270 182.915 ;
        RECT 214.440 182.775 214.615 183.105 ;
        RECT 215.320 183.035 215.490 184.205 ;
        RECT 216.405 184.115 217.055 184.285 ;
        RECT 216.120 183.555 216.575 183.725 ;
        RECT 215.900 183.375 216.310 183.385 ;
        RECT 215.900 183.215 216.315 183.375 ;
        RECT 216.885 183.335 217.055 184.115 ;
        RECT 216.140 183.045 216.315 183.215 ;
        RECT 216.485 183.165 217.055 183.335 ;
        RECT 214.960 182.865 215.490 183.035 ;
        RECT 215.660 182.875 215.830 183.035 ;
        RECT 216.485 182.875 216.655 183.165 ;
        RECT 214.960 182.705 215.130 182.865 ;
        RECT 215.660 182.705 216.655 182.875 ;
        RECT 216.825 182.535 216.995 182.995 ;
        RECT 217.245 182.705 217.505 184.915 ;
        RECT 217.765 184.155 217.935 184.915 ;
        RECT 218.115 184.325 218.445 185.085 ;
        RECT 217.765 183.985 218.430 184.155 ;
        RECT 218.615 184.010 218.885 184.915 ;
        RECT 220.065 184.415 220.235 184.915 ;
        RECT 220.405 184.705 220.735 185.085 ;
        RECT 220.905 184.745 222.435 184.915 ;
        RECT 220.905 184.585 221.075 184.745 ;
        RECT 221.425 184.415 221.595 184.575 ;
        RECT 220.065 184.245 221.595 184.415 ;
        RECT 221.765 184.405 222.095 184.575 ;
        RECT 221.765 184.075 221.935 184.405 ;
        RECT 222.265 184.245 222.435 184.745 ;
        RECT 222.605 184.075 222.955 184.915 ;
        RECT 223.125 184.705 223.455 185.085 ;
        RECT 223.715 184.745 224.725 184.915 ;
        RECT 218.260 183.840 218.430 183.985 ;
        RECT 217.695 183.435 218.025 183.805 ;
        RECT 218.260 183.510 218.545 183.840 ;
        RECT 218.260 183.255 218.430 183.510 ;
        RECT 217.765 183.085 218.430 183.255 ;
        RECT 218.715 183.210 218.885 184.010 ;
        RECT 220.035 183.895 220.385 184.065 ;
        RECT 220.040 183.445 220.385 183.895 ;
        RECT 220.695 183.445 221.130 184.065 ;
        RECT 221.300 183.905 221.935 184.075 ;
        RECT 221.300 183.385 221.470 183.905 ;
        RECT 222.150 183.845 222.955 184.075 ;
        RECT 222.150 183.735 222.510 183.845 ;
        RECT 221.970 183.555 222.510 183.735 ;
        RECT 217.765 182.705 217.935 183.085 ;
        RECT 218.115 182.535 218.445 182.915 ;
        RECT 218.625 182.705 218.885 183.210 ;
        RECT 220.065 183.085 221.075 183.255 ;
        RECT 220.065 182.710 220.235 183.085 ;
        RECT 220.405 182.535 220.735 182.915 ;
        RECT 220.905 182.875 221.075 183.085 ;
        RECT 221.300 183.215 221.590 183.385 ;
        RECT 221.300 183.045 221.640 183.215 ;
        RECT 221.810 182.875 221.980 183.210 ;
        RECT 222.150 182.880 222.510 183.555 ;
        RECT 223.155 183.445 223.455 184.445 ;
        RECT 223.715 184.235 223.885 184.745 ;
        RECT 224.055 184.065 224.385 184.575 ;
        RECT 224.555 184.535 224.725 184.745 ;
        RECT 224.950 184.705 225.280 185.085 ;
        RECT 225.450 184.535 225.620 184.915 ;
        RECT 225.870 184.705 226.220 185.085 ;
        RECT 226.390 184.585 226.575 184.915 ;
        RECT 224.555 184.365 225.620 184.535 ;
        RECT 224.690 184.065 224.935 184.125 ;
        RECT 223.625 183.895 224.385 184.065 ;
        RECT 224.635 183.895 224.935 184.065 ;
        RECT 223.625 183.370 223.795 183.895 ;
        RECT 224.180 183.715 224.350 183.725 ;
        RECT 223.965 183.555 224.350 183.715 ;
        RECT 223.965 183.545 224.295 183.555 ;
        RECT 224.690 183.505 224.935 183.895 ;
        RECT 225.140 184.065 225.470 184.125 ;
        RECT 225.140 183.895 225.495 184.065 ;
        RECT 225.140 183.505 225.470 183.895 ;
        RECT 225.945 183.445 226.235 184.125 ;
        RECT 226.405 183.725 226.575 184.585 ;
        RECT 226.870 184.585 227.080 184.915 ;
        RECT 227.250 184.745 228.535 184.915 ;
        RECT 227.250 184.705 227.580 184.745 ;
        RECT 226.405 183.555 226.695 183.725 ;
        RECT 223.625 183.295 223.940 183.370 ;
        RECT 220.905 182.705 221.980 182.875 ;
        RECT 222.690 182.535 222.980 183.255 ;
        RECT 223.270 182.875 223.440 183.245 ;
        RECT 223.610 183.045 223.940 183.295 ;
        RECT 224.110 183.335 224.280 183.375 ;
        RECT 224.110 183.165 225.630 183.335 ;
        RECT 224.110 183.045 224.280 183.165 ;
        RECT 224.515 182.875 224.870 182.915 ;
        RECT 223.270 182.705 224.870 182.875 ;
        RECT 225.040 182.535 225.210 182.995 ;
        RECT 225.385 182.745 225.630 183.165 ;
        RECT 226.405 183.105 226.575 183.555 ;
        RECT 226.870 183.385 227.040 184.585 ;
        RECT 227.735 184.435 228.065 184.575 ;
        RECT 227.280 184.205 228.065 184.435 ;
        RECT 228.365 184.285 228.535 184.745 ;
        RECT 228.705 184.705 229.035 185.085 ;
        RECT 226.870 183.215 227.110 183.385 ;
        RECT 225.900 182.535 226.230 182.915 ;
        RECT 226.400 182.775 226.575 183.105 ;
        RECT 227.280 183.035 227.450 184.205 ;
        RECT 228.365 184.115 229.015 184.285 ;
        RECT 228.080 183.555 228.535 183.725 ;
        RECT 227.860 183.375 228.270 183.385 ;
        RECT 227.860 183.215 228.275 183.375 ;
        RECT 228.845 183.335 229.015 184.115 ;
        RECT 228.100 183.045 228.275 183.215 ;
        RECT 228.445 183.165 229.015 183.335 ;
        RECT 226.920 182.865 227.450 183.035 ;
        RECT 227.620 182.875 227.790 183.035 ;
        RECT 228.445 182.875 228.615 183.165 ;
        RECT 226.920 182.705 227.090 182.865 ;
        RECT 227.620 182.705 228.615 182.875 ;
        RECT 228.785 182.535 228.955 182.995 ;
        RECT 229.205 182.705 229.465 184.915 ;
        RECT 229.635 183.920 229.925 185.085 ;
        RECT 230.095 184.010 230.365 184.915 ;
        RECT 230.535 184.325 230.865 185.085 ;
        RECT 231.045 184.155 231.215 184.915 ;
        RECT 229.635 182.535 229.925 183.260 ;
        RECT 230.095 183.210 230.265 184.010 ;
        RECT 230.550 183.985 231.215 184.155 ;
        RECT 231.475 184.010 231.745 184.915 ;
        RECT 231.915 184.325 232.245 185.085 ;
        RECT 232.425 184.155 232.595 184.915 ;
        RECT 230.550 183.840 230.720 183.985 ;
        RECT 230.435 183.510 230.720 183.840 ;
        RECT 230.550 183.255 230.720 183.510 ;
        RECT 230.955 183.435 231.285 183.805 ;
        RECT 230.095 182.705 230.355 183.210 ;
        RECT 230.550 183.085 231.215 183.255 ;
        RECT 230.535 182.535 230.865 182.915 ;
        RECT 231.045 182.705 231.215 183.085 ;
        RECT 231.475 183.210 231.645 184.010 ;
        RECT 231.930 183.985 232.595 184.155 ;
        RECT 232.855 184.010 233.125 184.915 ;
        RECT 233.295 184.325 233.625 185.085 ;
        RECT 233.805 184.155 233.975 184.915 ;
        RECT 231.930 183.840 232.100 183.985 ;
        RECT 231.815 183.510 232.100 183.840 ;
        RECT 231.930 183.255 232.100 183.510 ;
        RECT 232.335 183.435 232.665 183.805 ;
        RECT 231.475 182.705 231.735 183.210 ;
        RECT 231.930 183.085 232.595 183.255 ;
        RECT 231.915 182.535 232.245 182.915 ;
        RECT 232.425 182.705 232.595 183.085 ;
        RECT 232.855 183.210 233.025 184.010 ;
        RECT 233.310 183.985 233.975 184.155 ;
        RECT 234.235 184.010 234.505 184.915 ;
        RECT 234.675 184.325 235.005 185.085 ;
        RECT 235.185 184.155 235.355 184.915 ;
        RECT 233.310 183.840 233.480 183.985 ;
        RECT 233.195 183.510 233.480 183.840 ;
        RECT 233.310 183.255 233.480 183.510 ;
        RECT 233.715 183.435 234.045 183.805 ;
        RECT 232.855 182.705 233.115 183.210 ;
        RECT 233.310 183.085 233.975 183.255 ;
        RECT 233.295 182.535 233.625 182.915 ;
        RECT 233.805 182.705 233.975 183.085 ;
        RECT 234.235 183.210 234.405 184.010 ;
        RECT 234.690 183.985 235.355 184.155 ;
        RECT 235.615 184.010 235.885 184.915 ;
        RECT 236.055 184.325 236.385 185.085 ;
        RECT 236.565 184.155 236.735 184.915 ;
        RECT 234.690 183.840 234.860 183.985 ;
        RECT 234.575 183.510 234.860 183.840 ;
        RECT 234.690 183.255 234.860 183.510 ;
        RECT 235.095 183.435 235.425 183.805 ;
        RECT 234.235 182.705 234.495 183.210 ;
        RECT 234.690 183.085 235.355 183.255 ;
        RECT 234.675 182.535 235.005 182.915 ;
        RECT 235.185 182.705 235.355 183.085 ;
        RECT 235.615 183.210 235.785 184.010 ;
        RECT 236.070 183.985 236.735 184.155 ;
        RECT 237.915 183.995 239.125 185.085 ;
        RECT 236.070 183.840 236.240 183.985 ;
        RECT 235.955 183.510 236.240 183.840 ;
        RECT 236.070 183.255 236.240 183.510 ;
        RECT 236.475 183.435 236.805 183.805 ;
        RECT 237.915 183.455 238.435 183.995 ;
        RECT 238.605 183.285 239.125 183.825 ;
        RECT 235.615 182.705 235.875 183.210 ;
        RECT 236.070 183.085 236.735 183.255 ;
        RECT 236.055 182.535 236.385 182.915 ;
        RECT 236.565 182.705 236.735 183.085 ;
        RECT 237.915 182.535 239.125 183.285 ;
        RECT 165.150 182.365 239.210 182.535 ;
        RECT 165.235 181.615 166.445 182.365 ;
        RECT 166.615 181.865 166.875 182.195 ;
        RECT 167.085 181.885 167.360 182.365 ;
        RECT 165.235 181.075 165.755 181.615 ;
        RECT 102.225 180.620 155.700 181.020 ;
        RECT 165.925 180.905 166.445 181.445 ;
        RECT 62.895 180.305 99.045 180.475 ;
        RECT 9.330 178.450 52.060 178.620 ;
        RECT 9.330 168.690 9.500 178.450 ;
        RECT 10.230 177.760 12.230 177.930 ;
        RECT 12.520 177.760 14.520 177.930 ;
        RECT 14.810 177.760 16.810 177.930 ;
        RECT 17.100 177.760 19.100 177.930 ;
        RECT 19.390 177.760 21.390 177.930 ;
        RECT 21.680 177.760 23.680 177.930 ;
        RECT 23.970 177.760 25.970 177.930 ;
        RECT 26.260 177.760 28.260 177.930 ;
        RECT 28.550 177.760 30.550 177.930 ;
        RECT 30.840 177.760 32.840 177.930 ;
        RECT 33.130 177.760 35.130 177.930 ;
        RECT 35.420 177.760 37.420 177.930 ;
        RECT 37.710 177.760 39.710 177.930 ;
        RECT 40.000 177.760 42.000 177.930 ;
        RECT 42.290 177.760 44.290 177.930 ;
        RECT 44.580 177.760 46.580 177.930 ;
        RECT 46.870 177.760 48.870 177.930 ;
        RECT 49.160 177.760 51.160 177.930 ;
        RECT 10.000 169.550 10.170 177.590 ;
        RECT 12.290 169.550 12.460 177.590 ;
        RECT 14.580 169.550 14.750 177.590 ;
        RECT 16.870 169.550 17.040 177.590 ;
        RECT 19.160 169.550 19.330 177.590 ;
        RECT 21.450 169.550 21.620 177.590 ;
        RECT 23.740 169.550 23.910 177.590 ;
        RECT 26.030 169.550 26.200 177.590 ;
        RECT 28.320 169.550 28.490 177.590 ;
        RECT 30.610 169.550 30.780 177.590 ;
        RECT 32.900 169.550 33.070 177.590 ;
        RECT 35.190 169.550 35.360 177.590 ;
        RECT 37.480 169.550 37.650 177.590 ;
        RECT 39.770 169.550 39.940 177.590 ;
        RECT 42.060 169.550 42.230 177.590 ;
        RECT 44.350 169.550 44.520 177.590 ;
        RECT 46.640 169.550 46.810 177.590 ;
        RECT 48.930 169.550 49.100 177.590 ;
        RECT 51.220 169.550 51.390 177.590 ;
        RECT 10.230 169.210 12.230 169.380 ;
        RECT 12.520 169.210 14.520 169.380 ;
        RECT 14.810 169.210 16.810 169.380 ;
        RECT 17.100 169.210 19.100 169.380 ;
        RECT 19.390 169.210 21.390 169.380 ;
        RECT 21.680 169.210 23.680 169.380 ;
        RECT 23.970 169.210 25.970 169.380 ;
        RECT 26.260 169.210 28.260 169.380 ;
        RECT 28.550 169.210 30.550 169.380 ;
        RECT 30.840 169.210 32.840 169.380 ;
        RECT 33.130 169.210 35.130 169.380 ;
        RECT 35.420 169.210 37.420 169.380 ;
        RECT 37.710 169.210 39.710 169.380 ;
        RECT 40.000 169.210 42.000 169.380 ;
        RECT 42.290 169.210 44.290 169.380 ;
        RECT 44.580 169.210 46.580 169.380 ;
        RECT 46.870 169.210 48.870 169.380 ;
        RECT 49.160 169.210 51.160 169.380 ;
        RECT 51.890 168.690 52.060 178.450 ;
        RECT 62.895 177.455 63.425 180.305 ;
        RECT 64.155 179.615 80.155 179.785 ;
        RECT 63.925 178.360 64.095 179.400 ;
        RECT 80.215 178.360 80.385 179.400 ;
        RECT 64.155 177.975 80.155 178.145 ;
        RECT 80.885 177.455 81.055 180.305 ;
        RECT 81.785 179.615 97.785 179.785 ;
        RECT 81.555 178.360 81.725 179.400 ;
        RECT 97.845 178.360 98.015 179.400 ;
        RECT 81.785 177.975 97.785 178.145 ;
        RECT 98.515 177.455 99.045 180.305 ;
        RECT 62.895 177.285 99.045 177.455 ;
        RECT 62.895 174.435 63.425 177.285 ;
        RECT 64.155 176.595 80.155 176.765 ;
        RECT 63.925 175.340 64.095 176.380 ;
        RECT 80.215 175.340 80.385 176.380 ;
        RECT 64.155 174.955 80.155 175.125 ;
        RECT 80.885 174.435 81.055 177.285 ;
        RECT 81.785 176.595 97.785 176.765 ;
        RECT 81.555 175.340 81.725 176.380 ;
        RECT 97.845 175.340 98.015 176.380 ;
        RECT 81.785 174.955 97.785 175.125 ;
        RECT 98.515 174.435 99.045 177.285 ;
        RECT 62.895 174.265 99.045 174.435 ;
        RECT 62.895 171.415 63.425 174.265 ;
        RECT 63.925 173.575 80.385 173.745 ;
        RECT 63.925 172.105 64.155 173.575 ;
        RECT 80.155 172.105 80.385 173.575 ;
        RECT 63.925 171.935 80.385 172.105 ;
        RECT 80.885 171.415 81.055 174.265 ;
        RECT 81.555 173.575 98.015 173.745 ;
        RECT 81.555 172.105 81.785 173.575 ;
        RECT 97.785 172.105 98.015 173.575 ;
        RECT 81.555 171.935 98.015 172.105 ;
        RECT 98.515 171.415 99.045 174.265 ;
        RECT 113.860 176.355 151.710 176.885 ;
        RECT 62.895 170.885 99.045 171.415 ;
        RECT 102.740 172.330 110.970 172.500 ;
        RECT 9.330 168.520 52.060 168.690 ;
        RECT 9.330 167.860 51.780 168.030 ;
        RECT 9.330 158.100 9.500 167.860 ;
        RECT 10.290 167.170 12.290 167.340 ;
        RECT 12.580 167.170 14.580 167.340 ;
        RECT 10.060 158.960 10.230 167.000 ;
        RECT 12.350 158.960 12.520 167.000 ;
        RECT 14.640 158.960 14.810 167.000 ;
        RECT 10.290 158.620 12.290 158.790 ;
        RECT 12.580 158.620 14.580 158.790 ;
        RECT 15.370 158.100 15.540 167.860 ;
        RECT 16.330 167.170 18.330 167.340 ;
        RECT 18.620 167.170 20.620 167.340 ;
        RECT 16.100 158.960 16.270 167.000 ;
        RECT 18.390 158.960 18.560 167.000 ;
        RECT 20.680 158.960 20.850 167.000 ;
        RECT 16.330 158.620 18.330 158.790 ;
        RECT 18.620 158.620 20.620 158.790 ;
        RECT 21.410 158.100 21.580 167.860 ;
        RECT 22.370 167.170 24.370 167.340 ;
        RECT 24.660 167.170 26.660 167.340 ;
        RECT 22.140 158.960 22.310 167.000 ;
        RECT 24.430 158.960 24.600 167.000 ;
        RECT 26.720 158.960 26.890 167.000 ;
        RECT 22.370 158.620 24.370 158.790 ;
        RECT 24.660 158.620 26.660 158.790 ;
        RECT 27.450 158.100 27.620 167.860 ;
        RECT 28.410 167.170 30.410 167.340 ;
        RECT 30.700 167.170 32.700 167.340 ;
        RECT 28.180 158.960 28.350 167.000 ;
        RECT 30.470 158.960 30.640 167.000 ;
        RECT 32.760 158.960 32.930 167.000 ;
        RECT 28.410 158.620 30.410 158.790 ;
        RECT 30.700 158.620 32.700 158.790 ;
        RECT 33.490 158.100 33.660 167.860 ;
        RECT 34.450 167.170 36.450 167.340 ;
        RECT 36.740 167.170 38.740 167.340 ;
        RECT 34.220 158.960 34.390 167.000 ;
        RECT 36.510 158.960 36.680 167.000 ;
        RECT 38.800 158.960 38.970 167.000 ;
        RECT 34.450 158.620 36.450 158.790 ;
        RECT 36.740 158.620 38.740 158.790 ;
        RECT 39.530 158.100 39.700 167.860 ;
        RECT 40.490 167.170 42.490 167.340 ;
        RECT 42.780 167.170 44.780 167.340 ;
        RECT 40.260 158.960 40.430 167.000 ;
        RECT 42.550 158.960 42.720 167.000 ;
        RECT 44.840 158.960 45.010 167.000 ;
        RECT 40.490 158.620 42.490 158.790 ;
        RECT 42.780 158.620 44.780 158.790 ;
        RECT 45.570 158.100 45.740 167.860 ;
        RECT 46.530 167.170 48.530 167.340 ;
        RECT 48.820 167.170 50.820 167.340 ;
        RECT 46.300 158.960 46.470 167.000 ;
        RECT 48.590 158.960 48.760 167.000 ;
        RECT 50.880 158.960 51.050 167.000 ;
        RECT 46.530 158.620 48.530 158.790 ;
        RECT 48.820 158.620 50.820 158.790 ;
        RECT 51.610 158.100 51.780 167.860 ;
        RECT 9.330 157.930 51.780 158.100 ;
        RECT 9.330 148.170 9.500 157.930 ;
        RECT 10.290 157.240 12.290 157.410 ;
        RECT 12.580 157.240 14.580 157.410 ;
        RECT 10.060 149.030 10.230 157.070 ;
        RECT 12.350 149.030 12.520 157.070 ;
        RECT 14.640 149.030 14.810 157.070 ;
        RECT 10.290 148.690 12.290 148.860 ;
        RECT 12.580 148.690 14.580 148.860 ;
        RECT 15.370 148.170 15.540 157.930 ;
        RECT 16.330 157.240 18.330 157.410 ;
        RECT 18.620 157.240 20.620 157.410 ;
        RECT 16.100 149.030 16.270 157.070 ;
        RECT 18.390 149.030 18.560 157.070 ;
        RECT 20.680 149.030 20.850 157.070 ;
        RECT 16.330 148.690 18.330 148.860 ;
        RECT 18.620 148.690 20.620 148.860 ;
        RECT 21.410 148.170 21.580 157.930 ;
        RECT 22.370 157.240 24.370 157.410 ;
        RECT 24.660 157.240 26.660 157.410 ;
        RECT 22.140 149.030 22.310 157.070 ;
        RECT 24.430 149.030 24.600 157.070 ;
        RECT 26.720 149.030 26.890 157.070 ;
        RECT 22.370 148.690 24.370 148.860 ;
        RECT 24.660 148.690 26.660 148.860 ;
        RECT 27.450 148.170 27.620 157.930 ;
        RECT 28.410 157.240 30.410 157.410 ;
        RECT 30.700 157.240 32.700 157.410 ;
        RECT 28.180 149.030 28.350 157.070 ;
        RECT 30.470 149.030 30.640 157.070 ;
        RECT 32.760 149.030 32.930 157.070 ;
        RECT 28.410 148.690 30.410 148.860 ;
        RECT 30.700 148.690 32.700 148.860 ;
        RECT 33.490 148.170 33.660 157.930 ;
        RECT 34.450 157.240 36.450 157.410 ;
        RECT 36.740 157.240 38.740 157.410 ;
        RECT 34.220 149.030 34.390 157.070 ;
        RECT 36.510 149.030 36.680 157.070 ;
        RECT 38.800 149.030 38.970 157.070 ;
        RECT 34.450 148.690 36.450 148.860 ;
        RECT 36.740 148.690 38.740 148.860 ;
        RECT 39.530 148.170 39.700 157.930 ;
        RECT 40.490 157.240 42.490 157.410 ;
        RECT 42.780 157.240 44.780 157.410 ;
        RECT 40.260 149.030 40.430 157.070 ;
        RECT 42.550 149.030 42.720 157.070 ;
        RECT 44.840 149.030 45.010 157.070 ;
        RECT 40.490 148.690 42.490 148.860 ;
        RECT 42.780 148.690 44.780 148.860 ;
        RECT 45.570 148.170 45.740 157.930 ;
        RECT 46.530 157.240 48.530 157.410 ;
        RECT 48.820 157.240 50.820 157.410 ;
        RECT 46.300 149.030 46.470 157.070 ;
        RECT 48.590 149.030 48.760 157.070 ;
        RECT 50.880 149.030 51.050 157.070 ;
        RECT 46.530 148.690 48.530 148.860 ;
        RECT 48.820 148.690 50.820 148.860 ;
        RECT 51.610 148.170 51.780 157.930 ;
        RECT 9.330 148.000 51.780 148.170 ;
        RECT 64.100 166.025 96.940 166.425 ;
        RECT 23.195 143.155 58.705 143.745 ;
        RECT 23.195 140.745 23.785 143.155 ;
        RECT 24.515 142.465 32.515 142.635 ;
        RECT 32.805 142.465 40.805 142.635 ;
        RECT 41.095 142.465 49.095 142.635 ;
        RECT 49.385 142.465 57.385 142.635 ;
        RECT 24.285 141.255 24.455 142.295 ;
        RECT 32.575 141.255 32.745 142.295 ;
        RECT 40.865 141.255 41.035 142.295 ;
        RECT 49.155 141.255 49.325 142.295 ;
        RECT 57.445 141.255 57.615 142.295 ;
        RECT 24.515 140.915 32.515 141.085 ;
        RECT 32.805 140.915 40.805 141.085 ;
        RECT 41.095 140.915 49.095 141.085 ;
        RECT 49.385 140.915 57.385 141.085 ;
        RECT 23.195 139.705 24.455 140.745 ;
        RECT 32.575 139.705 32.745 140.745 ;
        RECT 40.865 139.705 41.035 140.745 ;
        RECT 49.155 139.705 49.325 140.745 ;
        RECT 57.445 139.705 57.615 140.745 ;
        RECT 23.195 139.195 23.785 139.705 ;
        RECT 24.515 139.365 32.515 139.535 ;
        RECT 32.805 139.365 40.805 139.535 ;
        RECT 41.095 139.365 49.095 139.535 ;
        RECT 49.385 139.365 57.385 139.535 ;
        RECT 9.430 137.955 20.720 138.485 ;
        RECT 9.430 135.195 9.960 137.955 ;
        RECT 10.995 137.265 11.995 137.435 ;
        RECT 10.765 136.055 10.935 137.095 ;
        RECT 12.055 136.055 12.225 137.095 ;
        RECT 13.030 135.195 13.200 137.955 ;
        RECT 13.930 137.265 14.930 137.435 ;
        RECT 15.220 137.265 16.220 137.435 ;
        RECT 13.700 136.055 13.870 137.095 ;
        RECT 14.990 136.055 15.160 137.095 ;
        RECT 16.280 136.055 16.450 137.095 ;
        RECT 16.950 135.195 17.120 137.955 ;
        RECT 18.155 137.265 19.155 137.435 ;
        RECT 17.925 136.055 18.095 137.095 ;
        RECT 19.215 136.055 19.385 137.095 ;
        RECT 20.190 135.195 20.720 137.955 ;
        RECT 9.430 134.665 20.720 135.195 ;
        RECT 23.195 138.155 24.455 139.195 ;
        RECT 32.575 138.155 32.745 139.195 ;
        RECT 40.865 138.155 41.035 139.195 ;
        RECT 49.155 138.155 49.325 139.195 ;
        RECT 57.445 138.155 57.615 139.195 ;
        RECT 23.195 135.745 23.785 138.155 ;
        RECT 24.515 137.815 32.515 137.985 ;
        RECT 32.805 137.815 40.805 137.985 ;
        RECT 41.095 137.815 49.095 137.985 ;
        RECT 49.385 137.815 57.385 137.985 ;
        RECT 24.285 136.605 24.455 137.645 ;
        RECT 32.575 136.605 32.745 137.645 ;
        RECT 40.865 136.605 41.035 137.645 ;
        RECT 49.155 136.605 49.325 137.645 ;
        RECT 57.445 136.605 57.615 137.645 ;
        RECT 24.515 136.265 32.515 136.435 ;
        RECT 32.805 136.265 40.805 136.435 ;
        RECT 41.095 136.265 49.095 136.435 ;
        RECT 49.385 136.265 57.385 136.435 ;
        RECT 58.115 135.745 58.705 143.155 ;
        RECT 23.195 135.155 58.705 135.745 ;
        RECT 64.100 133.985 64.500 166.025 ;
        RECT 69.635 160.720 91.405 160.890 ;
        RECT 69.635 139.290 69.805 160.720 ;
        RECT 71.220 158.800 89.820 159.305 ;
        RECT 71.220 156.090 71.725 158.800 ;
        RECT 72.035 158.130 74.125 158.490 ;
        RECT 72.035 156.760 72.395 158.130 ;
        RECT 72.685 157.050 73.475 157.840 ;
        RECT 73.765 156.760 74.125 158.130 ;
        RECT 72.035 156.400 74.125 156.760 ;
        RECT 74.435 156.090 75.445 158.800 ;
        RECT 75.755 158.130 77.845 158.490 ;
        RECT 75.755 156.760 76.115 158.130 ;
        RECT 76.405 157.050 77.195 157.840 ;
        RECT 77.485 156.760 77.845 158.130 ;
        RECT 75.755 156.400 77.845 156.760 ;
        RECT 78.155 156.090 79.165 158.800 ;
        RECT 79.475 158.130 81.565 158.490 ;
        RECT 79.475 156.760 79.835 158.130 ;
        RECT 80.125 157.050 80.915 157.840 ;
        RECT 81.205 156.760 81.565 158.130 ;
        RECT 79.475 156.400 81.565 156.760 ;
        RECT 81.875 156.090 82.885 158.800 ;
        RECT 83.195 158.130 85.285 158.490 ;
        RECT 83.195 156.760 83.555 158.130 ;
        RECT 83.845 157.050 84.635 157.840 ;
        RECT 84.925 156.760 85.285 158.130 ;
        RECT 83.195 156.400 85.285 156.760 ;
        RECT 85.595 156.090 86.605 158.800 ;
        RECT 86.915 158.130 89.005 158.490 ;
        RECT 86.915 156.760 87.275 158.130 ;
        RECT 87.565 157.050 88.355 157.840 ;
        RECT 88.645 156.760 89.005 158.130 ;
        RECT 86.915 156.400 89.005 156.760 ;
        RECT 89.315 156.090 89.820 158.800 ;
        RECT 71.220 155.080 89.820 156.090 ;
        RECT 71.220 152.370 71.725 155.080 ;
        RECT 72.035 154.410 74.125 154.770 ;
        RECT 72.035 153.040 72.395 154.410 ;
        RECT 72.685 153.330 73.475 154.120 ;
        RECT 73.765 153.040 74.125 154.410 ;
        RECT 72.035 152.680 74.125 153.040 ;
        RECT 74.435 152.370 75.445 155.080 ;
        RECT 75.755 154.410 77.845 154.770 ;
        RECT 75.755 153.040 76.115 154.410 ;
        RECT 76.405 153.330 77.195 154.120 ;
        RECT 77.485 153.040 77.845 154.410 ;
        RECT 75.755 152.680 77.845 153.040 ;
        RECT 78.155 152.370 79.165 155.080 ;
        RECT 79.475 154.410 81.565 154.770 ;
        RECT 79.475 153.040 79.835 154.410 ;
        RECT 80.125 153.330 80.915 154.120 ;
        RECT 81.205 153.040 81.565 154.410 ;
        RECT 79.475 152.680 81.565 153.040 ;
        RECT 81.875 152.370 82.885 155.080 ;
        RECT 83.195 154.410 85.285 154.770 ;
        RECT 83.195 153.040 83.555 154.410 ;
        RECT 83.845 153.330 84.635 154.120 ;
        RECT 84.925 153.040 85.285 154.410 ;
        RECT 83.195 152.680 85.285 153.040 ;
        RECT 85.595 152.370 86.605 155.080 ;
        RECT 86.915 154.410 89.005 154.770 ;
        RECT 86.915 153.040 87.275 154.410 ;
        RECT 87.565 153.330 88.355 154.120 ;
        RECT 88.645 153.040 89.005 154.410 ;
        RECT 86.915 152.680 89.005 153.040 ;
        RECT 89.315 152.370 89.820 155.080 ;
        RECT 71.220 151.360 89.820 152.370 ;
        RECT 71.220 148.650 71.725 151.360 ;
        RECT 72.035 150.690 74.125 151.050 ;
        RECT 72.035 149.320 72.395 150.690 ;
        RECT 72.685 149.610 73.475 150.400 ;
        RECT 73.765 149.320 74.125 150.690 ;
        RECT 72.035 148.960 74.125 149.320 ;
        RECT 74.435 148.650 75.445 151.360 ;
        RECT 75.755 150.690 77.845 151.050 ;
        RECT 75.755 149.320 76.115 150.690 ;
        RECT 76.405 149.610 77.195 150.400 ;
        RECT 77.485 149.320 77.845 150.690 ;
        RECT 75.755 148.960 77.845 149.320 ;
        RECT 78.155 148.650 79.165 151.360 ;
        RECT 79.475 150.690 81.565 151.050 ;
        RECT 79.475 149.320 79.835 150.690 ;
        RECT 80.125 149.610 80.915 150.400 ;
        RECT 81.205 149.320 81.565 150.690 ;
        RECT 79.475 148.960 81.565 149.320 ;
        RECT 81.875 148.650 82.885 151.360 ;
        RECT 83.195 150.690 85.285 151.050 ;
        RECT 83.195 149.320 83.555 150.690 ;
        RECT 83.845 149.610 84.635 150.400 ;
        RECT 84.925 149.320 85.285 150.690 ;
        RECT 83.195 148.960 85.285 149.320 ;
        RECT 85.595 148.650 86.605 151.360 ;
        RECT 86.915 150.690 89.005 151.050 ;
        RECT 86.915 149.320 87.275 150.690 ;
        RECT 87.565 149.610 88.355 150.400 ;
        RECT 88.645 149.320 89.005 150.690 ;
        RECT 86.915 148.960 89.005 149.320 ;
        RECT 89.315 148.650 89.820 151.360 ;
        RECT 71.220 147.640 89.820 148.650 ;
        RECT 71.220 144.930 71.725 147.640 ;
        RECT 72.035 146.970 74.125 147.330 ;
        RECT 72.035 145.600 72.395 146.970 ;
        RECT 72.685 145.890 73.475 146.680 ;
        RECT 73.765 145.600 74.125 146.970 ;
        RECT 72.035 145.240 74.125 145.600 ;
        RECT 74.435 144.930 75.445 147.640 ;
        RECT 75.755 146.970 77.845 147.330 ;
        RECT 75.755 145.600 76.115 146.970 ;
        RECT 76.405 145.890 77.195 146.680 ;
        RECT 77.485 145.600 77.845 146.970 ;
        RECT 75.755 145.240 77.845 145.600 ;
        RECT 78.155 144.930 79.165 147.640 ;
        RECT 79.475 146.970 81.565 147.330 ;
        RECT 79.475 145.600 79.835 146.970 ;
        RECT 80.125 145.890 80.915 146.680 ;
        RECT 81.205 145.600 81.565 146.970 ;
        RECT 79.475 145.240 81.565 145.600 ;
        RECT 81.875 144.930 82.885 147.640 ;
        RECT 83.195 146.970 85.285 147.330 ;
        RECT 83.195 145.600 83.555 146.970 ;
        RECT 83.845 145.890 84.635 146.680 ;
        RECT 84.925 145.600 85.285 146.970 ;
        RECT 83.195 145.240 85.285 145.600 ;
        RECT 85.595 144.930 86.605 147.640 ;
        RECT 86.915 146.970 89.005 147.330 ;
        RECT 86.915 145.600 87.275 146.970 ;
        RECT 87.565 145.890 88.355 146.680 ;
        RECT 88.645 145.600 89.005 146.970 ;
        RECT 86.915 145.240 89.005 145.600 ;
        RECT 89.315 144.930 89.820 147.640 ;
        RECT 71.220 143.920 89.820 144.930 ;
        RECT 71.220 141.210 71.725 143.920 ;
        RECT 72.035 143.250 74.125 143.610 ;
        RECT 72.035 141.880 72.395 143.250 ;
        RECT 72.685 142.170 73.475 142.960 ;
        RECT 73.765 141.880 74.125 143.250 ;
        RECT 72.035 141.520 74.125 141.880 ;
        RECT 74.435 141.210 75.445 143.920 ;
        RECT 75.755 143.250 77.845 143.610 ;
        RECT 75.755 141.880 76.115 143.250 ;
        RECT 76.405 142.170 77.195 142.960 ;
        RECT 77.485 141.880 77.845 143.250 ;
        RECT 75.755 141.520 77.845 141.880 ;
        RECT 78.155 141.210 79.165 143.920 ;
        RECT 79.475 143.250 81.565 143.610 ;
        RECT 79.475 141.880 79.835 143.250 ;
        RECT 80.125 142.170 80.915 142.960 ;
        RECT 81.205 141.880 81.565 143.250 ;
        RECT 79.475 141.520 81.565 141.880 ;
        RECT 81.875 141.210 82.885 143.920 ;
        RECT 83.195 143.250 85.285 143.610 ;
        RECT 83.195 141.880 83.555 143.250 ;
        RECT 83.845 142.170 84.635 142.960 ;
        RECT 84.925 141.880 85.285 143.250 ;
        RECT 83.195 141.520 85.285 141.880 ;
        RECT 85.595 141.210 86.605 143.920 ;
        RECT 86.915 143.250 89.005 143.610 ;
        RECT 86.915 141.880 87.275 143.250 ;
        RECT 87.565 142.170 88.355 142.960 ;
        RECT 88.645 141.880 89.005 143.250 ;
        RECT 86.915 141.520 89.005 141.880 ;
        RECT 89.315 141.210 89.820 143.920 ;
        RECT 71.220 140.705 89.820 141.210 ;
        RECT 91.235 139.290 91.405 160.720 ;
        RECT 69.635 139.120 91.405 139.290 ;
        RECT 96.540 133.985 96.940 166.025 ;
        RECT 102.740 162.570 102.910 172.330 ;
        RECT 103.695 171.640 104.695 171.810 ;
        RECT 104.985 171.640 105.985 171.810 ;
        RECT 103.465 163.430 103.635 171.470 ;
        RECT 104.755 163.430 104.925 171.470 ;
        RECT 106.045 163.430 106.215 171.470 ;
        RECT 103.695 163.090 104.695 163.260 ;
        RECT 104.985 163.090 105.985 163.260 ;
        RECT 106.770 162.570 106.940 172.330 ;
        RECT 107.725 171.640 108.725 171.810 ;
        RECT 109.015 171.640 110.015 171.810 ;
        RECT 107.495 163.430 107.665 171.470 ;
        RECT 108.785 163.430 108.955 171.470 ;
        RECT 110.075 163.430 110.245 171.470 ;
        RECT 107.725 163.090 108.725 163.260 ;
        RECT 109.015 163.090 110.015 163.260 ;
        RECT 110.800 162.570 110.970 172.330 ;
        RECT 113.860 166.595 114.390 176.355 ;
        RECT 115.180 175.665 115.680 175.835 ;
        RECT 115.970 175.665 116.470 175.835 ;
        RECT 116.760 175.665 117.260 175.835 ;
        RECT 117.550 175.665 118.050 175.835 ;
        RECT 114.950 167.455 115.120 175.495 ;
        RECT 115.740 167.455 115.910 175.495 ;
        RECT 116.530 167.455 116.700 175.495 ;
        RECT 117.320 167.455 117.490 175.495 ;
        RECT 118.110 167.455 118.280 175.495 ;
        RECT 115.180 167.115 115.680 167.285 ;
        RECT 115.970 167.115 116.470 167.285 ;
        RECT 116.760 167.115 117.260 167.285 ;
        RECT 117.550 167.115 118.050 167.285 ;
        RECT 118.840 166.595 119.010 176.355 ;
        RECT 119.800 175.665 120.300 175.835 ;
        RECT 120.590 175.665 121.090 175.835 ;
        RECT 121.380 175.665 121.880 175.835 ;
        RECT 122.170 175.665 122.670 175.835 ;
        RECT 119.570 167.455 119.740 175.495 ;
        RECT 120.360 167.455 120.530 175.495 ;
        RECT 121.150 167.455 121.320 175.495 ;
        RECT 121.940 167.455 122.110 175.495 ;
        RECT 122.730 167.455 122.900 175.495 ;
        RECT 119.800 167.115 120.300 167.285 ;
        RECT 120.590 167.115 121.090 167.285 ;
        RECT 121.380 167.115 121.880 167.285 ;
        RECT 122.170 167.115 122.670 167.285 ;
        RECT 123.460 166.595 123.630 176.355 ;
        RECT 124.420 175.665 124.920 175.835 ;
        RECT 125.210 175.665 125.710 175.835 ;
        RECT 126.000 175.665 126.500 175.835 ;
        RECT 126.790 175.665 127.290 175.835 ;
        RECT 124.190 167.455 124.360 175.495 ;
        RECT 124.980 167.455 125.150 175.495 ;
        RECT 125.770 167.455 125.940 175.495 ;
        RECT 126.560 167.455 126.730 175.495 ;
        RECT 127.350 167.455 127.520 175.495 ;
        RECT 124.420 167.115 124.920 167.285 ;
        RECT 125.210 167.115 125.710 167.285 ;
        RECT 126.000 167.115 126.500 167.285 ;
        RECT 126.790 167.115 127.290 167.285 ;
        RECT 128.080 166.595 128.250 176.355 ;
        RECT 129.040 175.665 129.540 175.835 ;
        RECT 129.830 175.665 130.330 175.835 ;
        RECT 130.620 175.665 131.120 175.835 ;
        RECT 131.410 175.665 131.910 175.835 ;
        RECT 128.810 167.455 128.980 175.495 ;
        RECT 129.600 167.455 129.770 175.495 ;
        RECT 130.390 167.455 130.560 175.495 ;
        RECT 131.180 167.455 131.350 175.495 ;
        RECT 131.970 167.455 132.140 175.495 ;
        RECT 129.040 167.115 129.540 167.285 ;
        RECT 129.830 167.115 130.330 167.285 ;
        RECT 130.620 167.115 131.120 167.285 ;
        RECT 131.410 167.115 131.910 167.285 ;
        RECT 132.700 166.595 132.870 176.355 ;
        RECT 133.660 175.665 134.160 175.835 ;
        RECT 134.450 175.665 134.950 175.835 ;
        RECT 135.240 175.665 135.740 175.835 ;
        RECT 136.030 175.665 136.530 175.835 ;
        RECT 133.430 167.455 133.600 175.495 ;
        RECT 134.220 167.455 134.390 175.495 ;
        RECT 135.010 167.455 135.180 175.495 ;
        RECT 135.800 167.455 135.970 175.495 ;
        RECT 136.590 167.455 136.760 175.495 ;
        RECT 133.660 167.115 134.160 167.285 ;
        RECT 134.450 167.115 134.950 167.285 ;
        RECT 135.240 167.115 135.740 167.285 ;
        RECT 136.030 167.115 136.530 167.285 ;
        RECT 137.320 166.595 137.490 176.355 ;
        RECT 138.280 175.665 138.780 175.835 ;
        RECT 139.070 175.665 139.570 175.835 ;
        RECT 139.860 175.665 140.360 175.835 ;
        RECT 140.650 175.665 141.150 175.835 ;
        RECT 138.050 167.455 138.220 175.495 ;
        RECT 138.840 167.455 139.010 175.495 ;
        RECT 139.630 167.455 139.800 175.495 ;
        RECT 140.420 167.455 140.590 175.495 ;
        RECT 141.210 167.455 141.380 175.495 ;
        RECT 138.280 167.115 138.780 167.285 ;
        RECT 139.070 167.115 139.570 167.285 ;
        RECT 139.860 167.115 140.360 167.285 ;
        RECT 140.650 167.115 141.150 167.285 ;
        RECT 141.940 166.595 142.110 176.355 ;
        RECT 142.900 175.665 143.400 175.835 ;
        RECT 143.690 175.665 144.190 175.835 ;
        RECT 144.480 175.665 144.980 175.835 ;
        RECT 145.270 175.665 145.770 175.835 ;
        RECT 142.670 167.455 142.840 175.495 ;
        RECT 143.460 167.455 143.630 175.495 ;
        RECT 144.250 167.455 144.420 175.495 ;
        RECT 145.040 167.455 145.210 175.495 ;
        RECT 145.830 167.455 146.000 175.495 ;
        RECT 142.900 167.115 143.400 167.285 ;
        RECT 143.690 167.115 144.190 167.285 ;
        RECT 144.480 167.115 144.980 167.285 ;
        RECT 145.270 167.115 145.770 167.285 ;
        RECT 146.560 166.595 146.730 176.355 ;
        RECT 147.520 175.665 148.020 175.835 ;
        RECT 148.310 175.665 148.810 175.835 ;
        RECT 149.100 175.665 149.600 175.835 ;
        RECT 149.890 175.665 150.390 175.835 ;
        RECT 147.290 167.455 147.460 175.495 ;
        RECT 148.080 167.455 148.250 175.495 ;
        RECT 148.870 167.455 149.040 175.495 ;
        RECT 149.660 167.455 149.830 175.495 ;
        RECT 150.450 167.455 150.620 175.495 ;
        RECT 147.520 167.115 148.020 167.285 ;
        RECT 148.310 167.115 148.810 167.285 ;
        RECT 149.100 167.115 149.600 167.285 ;
        RECT 149.890 167.115 150.390 167.285 ;
        RECT 151.180 166.595 151.710 176.355 ;
        RECT 113.860 166.065 151.710 166.595 ;
        RECT 102.740 162.400 110.970 162.570 ;
        RECT 102.740 158.640 102.910 162.400 ;
        RECT 103.465 159.500 103.635 161.540 ;
        RECT 104.755 159.500 104.925 161.540 ;
        RECT 106.045 159.500 106.215 161.540 ;
        RECT 103.695 159.160 104.695 159.330 ;
        RECT 104.985 159.160 105.985 159.330 ;
        RECT 106.770 158.640 106.940 162.400 ;
        RECT 107.495 159.500 107.665 161.540 ;
        RECT 108.785 159.500 108.955 161.540 ;
        RECT 110.075 159.500 110.245 161.540 ;
        RECT 107.725 159.160 108.725 159.330 ;
        RECT 109.015 159.160 110.015 159.330 ;
        RECT 110.800 158.640 110.970 162.400 ;
        RECT 102.740 158.470 110.970 158.640 ;
        RECT 116.015 157.500 149.445 158.030 ;
        RECT 102.740 155.775 110.970 155.945 ;
        RECT 102.740 151.925 102.910 155.775 ;
        RECT 103.695 155.085 104.695 155.255 ;
        RECT 104.985 155.085 105.985 155.255 ;
        RECT 103.465 152.830 103.635 154.870 ;
        RECT 104.755 152.830 104.925 154.870 ;
        RECT 106.045 152.830 106.215 154.870 ;
        RECT 106.770 151.925 106.940 155.775 ;
        RECT 107.725 155.085 108.725 155.255 ;
        RECT 109.015 155.085 110.015 155.255 ;
        RECT 107.495 152.830 107.665 154.870 ;
        RECT 108.785 152.830 108.955 154.870 ;
        RECT 110.075 152.830 110.245 154.870 ;
        RECT 110.800 151.925 110.970 155.775 ;
        RECT 102.740 151.755 110.970 151.925 ;
        RECT 102.740 141.905 102.910 151.755 ;
        RECT 103.695 151.065 104.695 151.235 ;
        RECT 104.985 151.065 105.985 151.235 ;
        RECT 103.465 142.810 103.635 150.850 ;
        RECT 104.755 142.810 104.925 150.850 ;
        RECT 106.045 142.810 106.215 150.850 ;
        RECT 103.695 142.425 104.695 142.595 ;
        RECT 104.985 142.425 105.985 142.595 ;
        RECT 106.770 141.905 106.940 151.755 ;
        RECT 107.725 151.065 108.725 151.235 ;
        RECT 109.015 151.065 110.015 151.235 ;
        RECT 107.495 142.810 107.665 150.850 ;
        RECT 108.785 142.810 108.955 150.850 ;
        RECT 110.075 142.810 110.245 150.850 ;
        RECT 107.725 142.425 108.725 142.595 ;
        RECT 109.015 142.425 110.015 142.595 ;
        RECT 110.800 141.905 110.970 151.755 ;
        RECT 102.740 141.735 110.970 141.905 ;
        RECT 116.015 140.250 116.545 157.500 ;
        RECT 117.130 156.135 119.290 156.825 ;
        RECT 117.130 154.965 119.290 155.655 ;
        RECT 117.130 153.795 119.290 154.485 ;
        RECT 117.130 152.625 119.290 153.315 ;
        RECT 117.130 151.455 119.290 152.145 ;
        RECT 117.130 150.285 119.290 150.975 ;
        RECT 117.130 149.115 119.290 149.805 ;
        RECT 117.130 147.945 119.290 148.635 ;
        RECT 117.130 146.775 119.290 147.465 ;
        RECT 117.130 145.605 119.290 146.295 ;
        RECT 117.130 144.435 119.290 145.125 ;
        RECT 117.130 143.265 119.290 143.955 ;
        RECT 117.130 142.095 119.290 142.785 ;
        RECT 117.130 140.925 119.290 141.615 ;
        RECT 119.595 140.250 122.075 157.500 ;
        RECT 122.380 156.135 124.540 156.825 ;
        RECT 125.060 156.135 127.220 156.825 ;
        RECT 122.380 154.965 124.540 155.655 ;
        RECT 125.060 154.965 127.220 155.655 ;
        RECT 122.380 153.795 124.540 154.485 ;
        RECT 125.060 153.795 127.220 154.485 ;
        RECT 122.380 152.625 124.540 153.315 ;
        RECT 125.060 152.625 127.220 153.315 ;
        RECT 122.380 151.455 124.540 152.145 ;
        RECT 125.060 151.455 127.220 152.145 ;
        RECT 122.380 150.285 124.540 150.975 ;
        RECT 125.060 150.285 127.220 150.975 ;
        RECT 122.380 149.115 124.540 149.805 ;
        RECT 125.060 149.115 127.220 149.805 ;
        RECT 122.380 147.945 124.540 148.635 ;
        RECT 125.060 147.945 127.220 148.635 ;
        RECT 122.380 146.775 124.540 147.465 ;
        RECT 125.060 146.775 127.220 147.465 ;
        RECT 122.380 145.605 124.540 146.295 ;
        RECT 125.060 145.605 127.220 146.295 ;
        RECT 122.380 144.435 124.540 145.125 ;
        RECT 125.060 144.435 127.220 145.125 ;
        RECT 122.380 143.265 124.540 143.955 ;
        RECT 125.060 143.265 127.220 143.955 ;
        RECT 122.380 142.095 124.540 142.785 ;
        RECT 125.060 142.095 127.220 142.785 ;
        RECT 122.380 140.925 124.540 141.615 ;
        RECT 125.060 140.925 127.220 141.615 ;
        RECT 127.525 140.250 130.005 157.500 ;
        RECT 130.310 156.135 132.470 156.825 ;
        RECT 132.990 156.135 135.150 156.825 ;
        RECT 130.310 154.965 132.470 155.655 ;
        RECT 132.990 154.965 135.150 155.655 ;
        RECT 130.310 153.795 132.470 154.485 ;
        RECT 132.990 153.795 135.150 154.485 ;
        RECT 130.310 152.625 132.470 153.315 ;
        RECT 132.990 152.625 135.150 153.315 ;
        RECT 130.310 151.455 132.470 152.145 ;
        RECT 132.990 151.455 135.150 152.145 ;
        RECT 130.310 150.285 132.470 150.975 ;
        RECT 132.990 150.285 135.150 150.975 ;
        RECT 130.310 149.115 132.470 149.805 ;
        RECT 132.990 149.115 135.150 149.805 ;
        RECT 130.310 147.945 132.470 148.635 ;
        RECT 132.990 147.945 135.150 148.635 ;
        RECT 130.310 146.775 132.470 147.465 ;
        RECT 132.990 146.775 135.150 147.465 ;
        RECT 130.310 145.605 132.470 146.295 ;
        RECT 132.990 145.605 135.150 146.295 ;
        RECT 130.310 144.435 132.470 145.125 ;
        RECT 132.990 144.435 135.150 145.125 ;
        RECT 130.310 143.265 132.470 143.955 ;
        RECT 132.990 143.265 135.150 143.955 ;
        RECT 130.310 142.095 132.470 142.785 ;
        RECT 132.990 142.095 135.150 142.785 ;
        RECT 130.310 140.925 132.470 141.615 ;
        RECT 132.990 140.925 135.150 141.615 ;
        RECT 135.455 140.250 137.935 157.500 ;
        RECT 138.240 156.135 140.400 156.825 ;
        RECT 140.920 156.135 143.080 156.825 ;
        RECT 138.240 154.965 140.400 155.655 ;
        RECT 140.920 154.965 143.080 155.655 ;
        RECT 138.240 153.795 140.400 154.485 ;
        RECT 140.920 153.795 143.080 154.485 ;
        RECT 138.240 152.625 140.400 153.315 ;
        RECT 140.920 152.625 143.080 153.315 ;
        RECT 138.240 151.455 140.400 152.145 ;
        RECT 140.920 151.455 143.080 152.145 ;
        RECT 138.240 150.285 140.400 150.975 ;
        RECT 140.920 150.285 143.080 150.975 ;
        RECT 138.240 149.115 140.400 149.805 ;
        RECT 140.920 149.115 143.080 149.805 ;
        RECT 138.240 147.945 140.400 148.635 ;
        RECT 140.920 147.945 143.080 148.635 ;
        RECT 138.240 146.775 140.400 147.465 ;
        RECT 140.920 146.775 143.080 147.465 ;
        RECT 138.240 145.605 140.400 146.295 ;
        RECT 140.920 145.605 143.080 146.295 ;
        RECT 138.240 144.435 140.400 145.125 ;
        RECT 140.920 144.435 143.080 145.125 ;
        RECT 138.240 143.265 140.400 143.955 ;
        RECT 140.920 143.265 143.080 143.955 ;
        RECT 138.240 142.095 140.400 142.785 ;
        RECT 140.920 142.095 143.080 142.785 ;
        RECT 138.240 140.925 140.400 141.615 ;
        RECT 140.920 140.925 143.080 141.615 ;
        RECT 143.385 140.250 145.865 157.500 ;
        RECT 146.170 156.135 148.330 156.825 ;
        RECT 146.170 154.965 148.330 155.655 ;
        RECT 146.170 153.795 148.330 154.485 ;
        RECT 146.170 152.625 148.330 153.315 ;
        RECT 146.170 151.455 148.330 152.145 ;
        RECT 146.170 150.285 148.330 150.975 ;
        RECT 146.170 149.115 148.330 149.805 ;
        RECT 146.170 147.945 148.330 148.635 ;
        RECT 146.170 146.775 148.330 147.465 ;
        RECT 146.170 145.605 148.330 146.295 ;
        RECT 146.170 144.435 148.330 145.125 ;
        RECT 146.170 143.265 148.330 143.955 ;
        RECT 146.170 142.095 148.330 142.785 ;
        RECT 146.170 140.925 148.330 141.615 ;
        RECT 148.915 140.250 149.445 157.500 ;
        RECT 116.015 139.720 149.445 140.250 ;
        RECT 64.100 133.585 96.940 133.985 ;
        RECT 138.110 134.130 145.930 134.660 ;
        RECT 138.110 130.280 138.640 134.130 ;
        RECT 139.465 133.440 140.465 133.610 ;
        RECT 140.755 133.440 141.755 133.610 ;
        RECT 139.235 131.185 139.405 133.225 ;
        RECT 140.525 131.185 140.695 133.225 ;
        RECT 141.815 131.185 141.985 133.225 ;
        RECT 142.580 130.280 142.750 134.130 ;
        RECT 143.345 131.185 143.515 133.225 ;
        RECT 144.635 131.185 144.805 133.225 ;
        RECT 143.575 130.800 144.575 130.970 ;
        RECT 145.400 130.280 145.930 134.130 ;
        RECT 138.110 129.750 145.930 130.280 ;
        RECT 138.110 128.410 145.930 128.940 ;
        RECT 138.110 124.650 138.640 128.410 ;
        RECT 139.235 125.510 139.405 127.550 ;
        RECT 140.525 125.510 140.695 127.550 ;
        RECT 141.815 125.510 141.985 127.550 ;
        RECT 139.465 125.170 140.465 125.340 ;
        RECT 140.755 125.170 141.755 125.340 ;
        RECT 142.580 124.650 142.750 128.410 ;
        RECT 143.575 127.720 144.575 127.890 ;
        RECT 143.345 125.510 143.515 127.550 ;
        RECT 144.635 125.510 144.805 127.550 ;
        RECT 145.400 124.650 145.930 128.410 ;
        RECT 10.055 123.725 70.145 124.255 ;
        RECT 10.055 113.875 10.585 123.725 ;
        RECT 11.315 123.035 13.315 123.205 ;
        RECT 13.605 123.035 15.605 123.205 ;
        RECT 11.085 114.780 11.255 122.820 ;
        RECT 13.375 114.780 13.545 122.820 ;
        RECT 15.665 114.780 15.835 122.820 ;
        RECT 11.315 114.395 13.315 114.565 ;
        RECT 13.605 114.395 15.605 114.565 ;
        RECT 16.335 113.875 16.505 123.725 ;
        RECT 17.235 123.035 19.235 123.205 ;
        RECT 19.525 123.035 21.525 123.205 ;
        RECT 17.005 114.780 17.175 122.820 ;
        RECT 19.295 114.780 19.465 122.820 ;
        RECT 21.585 114.780 21.755 122.820 ;
        RECT 17.235 114.395 19.235 114.565 ;
        RECT 19.525 114.395 21.525 114.565 ;
        RECT 22.255 113.875 22.425 123.725 ;
        RECT 23.155 123.035 25.155 123.205 ;
        RECT 25.445 123.035 27.445 123.205 ;
        RECT 22.925 114.780 23.095 122.820 ;
        RECT 25.215 114.780 25.385 122.820 ;
        RECT 27.505 114.780 27.675 122.820 ;
        RECT 23.155 114.395 25.155 114.565 ;
        RECT 25.445 114.395 27.445 114.565 ;
        RECT 28.175 113.875 28.345 123.725 ;
        RECT 29.075 123.035 31.075 123.205 ;
        RECT 31.365 123.035 33.365 123.205 ;
        RECT 28.845 114.780 29.015 122.820 ;
        RECT 31.135 114.780 31.305 122.820 ;
        RECT 33.425 114.780 33.595 122.820 ;
        RECT 29.075 114.395 31.075 114.565 ;
        RECT 31.365 114.395 33.365 114.565 ;
        RECT 34.095 113.875 34.265 123.725 ;
        RECT 34.995 123.035 36.995 123.205 ;
        RECT 37.285 123.035 39.285 123.205 ;
        RECT 34.765 114.780 34.935 122.820 ;
        RECT 37.055 114.780 37.225 122.820 ;
        RECT 39.345 114.780 39.515 122.820 ;
        RECT 34.995 114.395 36.995 114.565 ;
        RECT 37.285 114.395 39.285 114.565 ;
        RECT 40.015 113.875 40.185 123.725 ;
        RECT 40.915 123.035 42.915 123.205 ;
        RECT 43.205 123.035 45.205 123.205 ;
        RECT 40.685 114.780 40.855 122.820 ;
        RECT 42.975 114.780 43.145 122.820 ;
        RECT 45.265 114.780 45.435 122.820 ;
        RECT 40.915 114.395 42.915 114.565 ;
        RECT 43.205 114.395 45.205 114.565 ;
        RECT 45.935 113.875 46.105 123.725 ;
        RECT 46.835 123.035 48.835 123.205 ;
        RECT 49.125 123.035 51.125 123.205 ;
        RECT 46.605 114.780 46.775 122.820 ;
        RECT 48.895 114.780 49.065 122.820 ;
        RECT 51.185 114.780 51.355 122.820 ;
        RECT 46.835 114.395 48.835 114.565 ;
        RECT 49.125 114.395 51.125 114.565 ;
        RECT 51.855 113.875 52.025 123.725 ;
        RECT 52.755 123.035 54.755 123.205 ;
        RECT 55.045 123.035 57.045 123.205 ;
        RECT 52.525 114.780 52.695 122.820 ;
        RECT 54.815 114.780 54.985 122.820 ;
        RECT 57.105 114.780 57.275 122.820 ;
        RECT 52.755 114.395 54.755 114.565 ;
        RECT 55.045 114.395 57.045 114.565 ;
        RECT 57.775 113.875 57.945 123.725 ;
        RECT 58.675 123.035 60.675 123.205 ;
        RECT 60.965 123.035 62.965 123.205 ;
        RECT 58.445 114.780 58.615 122.820 ;
        RECT 60.735 114.780 60.905 122.820 ;
        RECT 63.025 114.780 63.195 122.820 ;
        RECT 58.675 114.395 60.675 114.565 ;
        RECT 60.965 114.395 62.965 114.565 ;
        RECT 63.695 113.875 63.865 123.725 ;
        RECT 64.595 123.035 66.595 123.205 ;
        RECT 66.885 123.035 68.885 123.205 ;
        RECT 64.365 114.780 64.535 122.820 ;
        RECT 66.655 114.780 66.825 122.820 ;
        RECT 68.945 114.780 69.115 122.820 ;
        RECT 64.595 114.395 66.595 114.565 ;
        RECT 66.885 114.395 68.885 114.565 ;
        RECT 69.615 113.875 70.145 123.725 ;
        RECT 10.055 113.705 70.145 113.875 ;
        RECT 10.055 103.855 10.585 113.705 ;
        RECT 11.315 113.015 13.315 113.185 ;
        RECT 13.605 113.015 15.605 113.185 ;
        RECT 11.085 104.760 11.255 112.800 ;
        RECT 13.375 104.760 13.545 112.800 ;
        RECT 15.665 104.760 15.835 112.800 ;
        RECT 11.315 104.375 13.315 104.545 ;
        RECT 13.605 104.375 15.605 104.545 ;
        RECT 16.335 103.855 16.505 113.705 ;
        RECT 17.235 113.015 19.235 113.185 ;
        RECT 19.525 113.015 21.525 113.185 ;
        RECT 17.005 104.760 17.175 112.800 ;
        RECT 19.295 104.760 19.465 112.800 ;
        RECT 21.585 104.760 21.755 112.800 ;
        RECT 17.235 104.375 19.235 104.545 ;
        RECT 19.525 104.375 21.525 104.545 ;
        RECT 22.255 103.855 22.425 113.705 ;
        RECT 23.155 113.015 25.155 113.185 ;
        RECT 25.445 113.015 27.445 113.185 ;
        RECT 22.925 104.760 23.095 112.800 ;
        RECT 25.215 104.760 25.385 112.800 ;
        RECT 27.505 104.760 27.675 112.800 ;
        RECT 23.155 104.375 25.155 104.545 ;
        RECT 25.445 104.375 27.445 104.545 ;
        RECT 28.175 103.855 28.345 113.705 ;
        RECT 29.075 113.015 31.075 113.185 ;
        RECT 31.365 113.015 33.365 113.185 ;
        RECT 28.845 104.760 29.015 112.800 ;
        RECT 31.135 104.760 31.305 112.800 ;
        RECT 33.425 104.760 33.595 112.800 ;
        RECT 29.075 104.375 31.075 104.545 ;
        RECT 31.365 104.375 33.365 104.545 ;
        RECT 34.095 103.855 34.265 113.705 ;
        RECT 34.995 113.015 36.995 113.185 ;
        RECT 37.285 113.015 39.285 113.185 ;
        RECT 34.765 104.760 34.935 112.800 ;
        RECT 37.055 104.760 37.225 112.800 ;
        RECT 39.345 104.760 39.515 112.800 ;
        RECT 34.995 104.375 36.995 104.545 ;
        RECT 37.285 104.375 39.285 104.545 ;
        RECT 40.015 103.855 40.185 113.705 ;
        RECT 40.915 113.015 42.915 113.185 ;
        RECT 43.205 113.015 45.205 113.185 ;
        RECT 40.685 104.760 40.855 112.800 ;
        RECT 42.975 104.760 43.145 112.800 ;
        RECT 45.265 104.760 45.435 112.800 ;
        RECT 40.915 104.375 42.915 104.545 ;
        RECT 43.205 104.375 45.205 104.545 ;
        RECT 45.935 103.855 46.105 113.705 ;
        RECT 46.835 113.015 48.835 113.185 ;
        RECT 49.125 113.015 51.125 113.185 ;
        RECT 46.605 104.760 46.775 112.800 ;
        RECT 48.895 104.760 49.065 112.800 ;
        RECT 51.185 104.760 51.355 112.800 ;
        RECT 46.835 104.375 48.835 104.545 ;
        RECT 49.125 104.375 51.125 104.545 ;
        RECT 51.855 103.855 52.025 113.705 ;
        RECT 52.755 113.015 54.755 113.185 ;
        RECT 55.045 113.015 57.045 113.185 ;
        RECT 52.525 104.760 52.695 112.800 ;
        RECT 54.815 104.760 54.985 112.800 ;
        RECT 57.105 104.760 57.275 112.800 ;
        RECT 52.755 104.375 54.755 104.545 ;
        RECT 55.045 104.375 57.045 104.545 ;
        RECT 57.775 103.855 57.945 113.705 ;
        RECT 58.675 113.015 60.675 113.185 ;
        RECT 60.965 113.015 62.965 113.185 ;
        RECT 58.445 104.760 58.615 112.800 ;
        RECT 60.735 104.760 60.905 112.800 ;
        RECT 63.025 104.760 63.195 112.800 ;
        RECT 58.675 104.375 60.675 104.545 ;
        RECT 60.965 104.375 62.965 104.545 ;
        RECT 63.695 103.855 63.865 113.705 ;
        RECT 64.595 113.015 66.595 113.185 ;
        RECT 66.885 113.015 68.885 113.185 ;
        RECT 64.365 104.760 64.535 112.800 ;
        RECT 66.655 104.760 66.825 112.800 ;
        RECT 68.945 104.760 69.115 112.800 ;
        RECT 64.595 104.375 66.595 104.545 ;
        RECT 66.885 104.375 68.885 104.545 ;
        RECT 69.615 103.855 70.145 113.705 ;
        RECT 10.055 103.325 70.145 103.855 ;
        RECT 71.805 123.725 114.135 124.255 ;
        RECT 138.110 124.120 145.930 124.650 ;
        RECT 71.805 113.875 72.335 123.725 ;
        RECT 72.835 122.820 77.585 123.725 ;
        RECT 72.835 114.780 73.005 122.820 ;
        RECT 75.125 114.780 75.295 122.820 ;
        RECT 77.415 114.780 77.585 122.820 ;
        RECT 73.065 114.395 75.065 114.565 ;
        RECT 75.355 114.395 77.355 114.565 ;
        RECT 78.085 113.875 78.255 123.725 ;
        RECT 78.985 123.035 80.985 123.205 ;
        RECT 81.275 123.035 83.275 123.205 ;
        RECT 78.755 114.780 78.925 122.820 ;
        RECT 81.045 114.780 81.215 122.820 ;
        RECT 83.335 114.780 83.505 122.820 ;
        RECT 78.985 114.395 80.985 114.565 ;
        RECT 81.275 114.395 83.275 114.565 ;
        RECT 84.005 113.875 84.175 123.725 ;
        RECT 84.905 123.035 86.905 123.205 ;
        RECT 87.195 123.035 89.195 123.205 ;
        RECT 84.675 114.780 84.845 122.820 ;
        RECT 86.965 114.780 87.135 122.820 ;
        RECT 89.255 114.780 89.425 122.820 ;
        RECT 84.905 114.395 86.905 114.565 ;
        RECT 87.195 114.395 89.195 114.565 ;
        RECT 89.925 113.875 90.095 123.725 ;
        RECT 90.825 123.035 92.825 123.205 ;
        RECT 93.115 123.035 95.115 123.205 ;
        RECT 90.595 114.780 90.765 122.820 ;
        RECT 92.885 114.780 93.055 122.820 ;
        RECT 95.175 114.780 95.345 122.820 ;
        RECT 90.825 114.395 92.825 114.565 ;
        RECT 93.115 114.395 95.115 114.565 ;
        RECT 95.845 113.875 96.015 123.725 ;
        RECT 96.745 123.035 98.745 123.205 ;
        RECT 99.035 123.035 101.035 123.205 ;
        RECT 96.515 114.780 96.685 122.820 ;
        RECT 98.805 114.780 98.975 122.820 ;
        RECT 101.095 114.780 101.265 122.820 ;
        RECT 96.745 114.395 98.745 114.565 ;
        RECT 99.035 114.395 101.035 114.565 ;
        RECT 101.765 113.875 101.935 123.725 ;
        RECT 102.665 123.035 104.665 123.205 ;
        RECT 104.955 123.035 106.955 123.205 ;
        RECT 102.435 114.780 102.605 122.820 ;
        RECT 104.725 114.780 104.895 122.820 ;
        RECT 107.015 114.780 107.185 122.820 ;
        RECT 102.665 114.395 104.665 114.565 ;
        RECT 104.955 114.395 106.955 114.565 ;
        RECT 107.685 113.875 107.855 123.725 ;
        RECT 108.355 122.820 113.105 123.725 ;
        RECT 108.355 114.780 108.525 122.820 ;
        RECT 110.645 114.780 110.815 122.820 ;
        RECT 112.935 114.780 113.105 122.820 ;
        RECT 108.585 114.395 110.585 114.565 ;
        RECT 110.875 114.395 112.875 114.565 ;
        RECT 113.605 113.875 114.135 123.725 ;
        RECT 71.805 113.705 114.135 113.875 ;
        RECT 71.805 103.855 72.335 113.705 ;
        RECT 73.065 113.015 75.065 113.185 ;
        RECT 75.355 113.015 77.355 113.185 ;
        RECT 72.835 104.760 73.005 112.800 ;
        RECT 75.125 104.760 75.295 112.800 ;
        RECT 77.415 104.760 77.585 112.800 ;
        RECT 72.835 103.855 77.585 104.760 ;
        RECT 78.085 103.855 78.255 113.705 ;
        RECT 78.985 113.015 80.985 113.185 ;
        RECT 81.275 113.015 83.275 113.185 ;
        RECT 78.755 104.760 78.925 112.800 ;
        RECT 81.045 104.760 81.215 112.800 ;
        RECT 83.335 104.760 83.505 112.800 ;
        RECT 78.985 104.375 80.985 104.545 ;
        RECT 81.275 104.375 83.275 104.545 ;
        RECT 84.005 103.855 84.175 113.705 ;
        RECT 84.905 113.015 86.905 113.185 ;
        RECT 87.195 113.015 89.195 113.185 ;
        RECT 84.675 104.760 84.845 112.800 ;
        RECT 86.965 104.760 87.135 112.800 ;
        RECT 89.255 104.760 89.425 112.800 ;
        RECT 84.905 104.375 86.905 104.545 ;
        RECT 87.195 104.375 89.195 104.545 ;
        RECT 89.925 103.855 90.095 113.705 ;
        RECT 90.825 113.015 92.825 113.185 ;
        RECT 93.115 113.015 95.115 113.185 ;
        RECT 90.595 104.760 90.765 112.800 ;
        RECT 92.885 104.760 93.055 112.800 ;
        RECT 95.175 104.760 95.345 112.800 ;
        RECT 90.825 104.375 92.825 104.545 ;
        RECT 93.115 104.375 95.115 104.545 ;
        RECT 95.845 103.855 96.015 113.705 ;
        RECT 96.745 113.015 98.745 113.185 ;
        RECT 99.035 113.015 101.035 113.185 ;
        RECT 96.515 104.760 96.685 112.800 ;
        RECT 98.805 104.760 98.975 112.800 ;
        RECT 101.095 104.760 101.265 112.800 ;
        RECT 96.745 104.375 98.745 104.545 ;
        RECT 99.035 104.375 101.035 104.545 ;
        RECT 101.765 103.855 101.935 113.705 ;
        RECT 102.665 113.015 104.665 113.185 ;
        RECT 104.955 113.015 106.955 113.185 ;
        RECT 102.435 104.760 102.605 112.800 ;
        RECT 104.725 104.760 104.895 112.800 ;
        RECT 107.015 104.760 107.185 112.800 ;
        RECT 102.665 104.375 104.665 104.545 ;
        RECT 104.955 104.375 106.955 104.545 ;
        RECT 107.685 103.855 107.855 113.705 ;
        RECT 108.585 113.015 110.585 113.185 ;
        RECT 110.875 113.015 112.875 113.185 ;
        RECT 108.355 104.760 108.525 112.800 ;
        RECT 110.645 104.760 110.815 112.800 ;
        RECT 112.935 104.760 113.105 112.800 ;
        RECT 108.355 103.855 113.105 104.760 ;
        RECT 113.605 103.855 114.135 113.705 ;
        RECT 71.805 103.325 114.135 103.855 ;
        RECT 115.935 122.945 128.905 123.475 ;
        RECT 115.935 113.485 116.465 122.945 ;
        RECT 117.370 122.275 118.410 122.445 ;
        RECT 116.985 114.215 117.155 122.215 ;
        RECT 118.625 114.215 118.795 122.215 ;
        RECT 117.370 113.985 118.410 114.155 ;
        RECT 119.315 113.485 119.485 122.945 ;
        RECT 120.390 122.275 121.430 122.445 ;
        RECT 120.005 114.215 120.175 122.215 ;
        RECT 121.645 114.215 121.815 122.215 ;
        RECT 120.390 113.985 121.430 114.155 ;
        RECT 122.335 113.485 122.505 122.945 ;
        RECT 123.410 122.275 124.450 122.445 ;
        RECT 123.025 114.215 123.195 122.215 ;
        RECT 124.665 114.215 124.835 122.215 ;
        RECT 123.410 113.985 124.450 114.155 ;
        RECT 125.355 113.485 125.525 122.945 ;
        RECT 126.430 122.275 127.470 122.445 ;
        RECT 126.045 114.215 126.215 122.215 ;
        RECT 127.685 114.215 127.855 122.215 ;
        RECT 126.430 113.985 127.470 114.155 ;
        RECT 128.375 113.485 128.905 122.945 ;
        RECT 115.935 113.315 128.905 113.485 ;
        RECT 115.935 103.855 116.465 113.315 ;
        RECT 117.370 112.645 118.410 112.815 ;
        RECT 116.985 104.585 117.155 112.585 ;
        RECT 118.625 104.585 118.795 112.585 ;
        RECT 117.370 104.355 118.410 104.525 ;
        RECT 119.315 103.855 119.485 113.315 ;
        RECT 120.390 112.645 121.430 112.815 ;
        RECT 120.005 104.585 120.175 112.585 ;
        RECT 121.645 104.585 121.815 112.585 ;
        RECT 120.390 104.355 121.430 104.525 ;
        RECT 122.335 103.855 122.505 113.315 ;
        RECT 123.410 112.645 124.450 112.815 ;
        RECT 123.025 104.585 123.195 112.585 ;
        RECT 124.665 104.585 124.835 112.585 ;
        RECT 123.410 104.355 124.450 104.525 ;
        RECT 125.355 103.855 125.525 113.315 ;
        RECT 126.430 112.645 127.470 112.815 ;
        RECT 126.045 104.585 126.215 112.585 ;
        RECT 127.685 104.585 127.855 112.585 ;
        RECT 126.430 104.355 127.470 104.525 ;
        RECT 128.375 103.855 128.905 113.315 ;
        RECT 115.935 103.325 128.905 103.855 ;
        RECT 135.150 104.785 149.540 108.660 ;
        RECT 10.055 102.145 128.905 102.675 ;
        RECT 10.055 92.295 10.585 102.145 ;
        RECT 11.315 101.455 13.315 101.625 ;
        RECT 13.605 101.455 15.605 101.625 ;
        RECT 15.895 101.455 17.895 101.625 ;
        RECT 18.185 101.455 20.185 101.625 ;
        RECT 20.475 101.455 22.475 101.625 ;
        RECT 22.765 101.455 24.765 101.625 ;
        RECT 25.055 101.455 27.055 101.625 ;
        RECT 27.345 101.455 29.345 101.625 ;
        RECT 11.085 93.200 11.255 101.240 ;
        RECT 13.375 93.200 13.545 101.240 ;
        RECT 15.665 93.200 15.835 101.240 ;
        RECT 17.955 93.200 18.125 101.240 ;
        RECT 20.245 93.200 20.415 101.240 ;
        RECT 22.535 93.200 22.705 101.240 ;
        RECT 24.825 93.200 24.995 101.240 ;
        RECT 27.115 93.200 27.285 101.240 ;
        RECT 29.405 93.200 29.575 101.240 ;
        RECT 11.315 92.815 13.315 92.985 ;
        RECT 13.605 92.815 15.605 92.985 ;
        RECT 15.895 92.815 17.895 92.985 ;
        RECT 18.185 92.815 20.185 92.985 ;
        RECT 20.475 92.815 22.475 92.985 ;
        RECT 22.765 92.815 24.765 92.985 ;
        RECT 25.055 92.815 27.055 92.985 ;
        RECT 27.345 92.815 29.345 92.985 ;
        RECT 30.075 92.295 30.245 102.145 ;
        RECT 30.975 101.455 32.975 101.625 ;
        RECT 33.265 101.455 35.265 101.625 ;
        RECT 35.555 101.455 37.555 101.625 ;
        RECT 37.845 101.455 39.845 101.625 ;
        RECT 40.135 101.455 42.135 101.625 ;
        RECT 42.425 101.455 44.425 101.625 ;
        RECT 44.715 101.455 46.715 101.625 ;
        RECT 47.005 101.455 49.005 101.625 ;
        RECT 30.745 93.200 30.915 101.240 ;
        RECT 33.035 93.200 33.205 101.240 ;
        RECT 35.325 93.200 35.495 101.240 ;
        RECT 37.615 93.200 37.785 101.240 ;
        RECT 39.905 93.200 40.075 101.240 ;
        RECT 42.195 93.200 42.365 101.240 ;
        RECT 44.485 93.200 44.655 101.240 ;
        RECT 46.775 93.200 46.945 101.240 ;
        RECT 49.065 93.200 49.235 101.240 ;
        RECT 30.975 92.815 32.975 92.985 ;
        RECT 33.265 92.815 35.265 92.985 ;
        RECT 35.555 92.815 37.555 92.985 ;
        RECT 37.845 92.815 39.845 92.985 ;
        RECT 40.135 92.815 42.135 92.985 ;
        RECT 42.425 92.815 44.425 92.985 ;
        RECT 44.715 92.815 46.715 92.985 ;
        RECT 47.005 92.815 49.005 92.985 ;
        RECT 49.735 92.295 49.905 102.145 ;
        RECT 50.635 101.455 52.635 101.625 ;
        RECT 52.925 101.455 54.925 101.625 ;
        RECT 55.215 101.455 57.215 101.625 ;
        RECT 57.505 101.455 59.505 101.625 ;
        RECT 59.795 101.455 61.795 101.625 ;
        RECT 62.085 101.455 64.085 101.625 ;
        RECT 64.375 101.455 66.375 101.625 ;
        RECT 66.665 101.455 68.665 101.625 ;
        RECT 50.405 93.200 50.575 101.240 ;
        RECT 52.695 93.200 52.865 101.240 ;
        RECT 54.985 93.200 55.155 101.240 ;
        RECT 57.275 93.200 57.445 101.240 ;
        RECT 59.565 93.200 59.735 101.240 ;
        RECT 61.855 93.200 62.025 101.240 ;
        RECT 64.145 93.200 64.315 101.240 ;
        RECT 66.435 93.200 66.605 101.240 ;
        RECT 68.725 93.200 68.895 101.240 ;
        RECT 50.635 92.815 52.635 92.985 ;
        RECT 52.925 92.815 54.925 92.985 ;
        RECT 55.215 92.815 57.215 92.985 ;
        RECT 57.505 92.815 59.505 92.985 ;
        RECT 59.795 92.815 61.795 92.985 ;
        RECT 62.085 92.815 64.085 92.985 ;
        RECT 64.375 92.815 66.375 92.985 ;
        RECT 66.665 92.815 68.665 92.985 ;
        RECT 69.395 92.295 69.565 102.145 ;
        RECT 70.295 101.455 72.295 101.625 ;
        RECT 72.585 101.455 74.585 101.625 ;
        RECT 74.875 101.455 76.875 101.625 ;
        RECT 77.165 101.455 79.165 101.625 ;
        RECT 79.455 101.455 81.455 101.625 ;
        RECT 81.745 101.455 83.745 101.625 ;
        RECT 84.035 101.455 86.035 101.625 ;
        RECT 86.325 101.455 88.325 101.625 ;
        RECT 70.065 93.200 70.235 101.240 ;
        RECT 72.355 93.200 72.525 101.240 ;
        RECT 74.645 93.200 74.815 101.240 ;
        RECT 76.935 93.200 77.105 101.240 ;
        RECT 79.225 93.200 79.395 101.240 ;
        RECT 81.515 93.200 81.685 101.240 ;
        RECT 83.805 93.200 83.975 101.240 ;
        RECT 86.095 93.200 86.265 101.240 ;
        RECT 88.385 93.200 88.555 101.240 ;
        RECT 70.295 92.815 72.295 92.985 ;
        RECT 72.585 92.815 74.585 92.985 ;
        RECT 74.875 92.815 76.875 92.985 ;
        RECT 77.165 92.815 79.165 92.985 ;
        RECT 79.455 92.815 81.455 92.985 ;
        RECT 81.745 92.815 83.745 92.985 ;
        RECT 84.035 92.815 86.035 92.985 ;
        RECT 86.325 92.815 88.325 92.985 ;
        RECT 89.055 92.295 89.225 102.145 ;
        RECT 89.955 101.455 91.955 101.625 ;
        RECT 92.245 101.455 94.245 101.625 ;
        RECT 94.535 101.455 96.535 101.625 ;
        RECT 96.825 101.455 98.825 101.625 ;
        RECT 99.115 101.455 101.115 101.625 ;
        RECT 101.405 101.455 103.405 101.625 ;
        RECT 103.695 101.455 105.695 101.625 ;
        RECT 105.985 101.455 107.985 101.625 ;
        RECT 89.725 93.200 89.895 101.240 ;
        RECT 92.015 93.200 92.185 101.240 ;
        RECT 94.305 93.200 94.475 101.240 ;
        RECT 96.595 93.200 96.765 101.240 ;
        RECT 98.885 93.200 99.055 101.240 ;
        RECT 101.175 93.200 101.345 101.240 ;
        RECT 103.465 93.200 103.635 101.240 ;
        RECT 105.755 93.200 105.925 101.240 ;
        RECT 108.045 93.200 108.215 101.240 ;
        RECT 89.955 92.815 91.955 92.985 ;
        RECT 92.245 92.815 94.245 92.985 ;
        RECT 94.535 92.815 96.535 92.985 ;
        RECT 96.825 92.815 98.825 92.985 ;
        RECT 99.115 92.815 101.115 92.985 ;
        RECT 101.405 92.815 103.405 92.985 ;
        RECT 103.695 92.815 105.695 92.985 ;
        RECT 105.985 92.815 107.985 92.985 ;
        RECT 108.715 92.295 108.885 102.145 ;
        RECT 109.615 101.455 111.615 101.625 ;
        RECT 111.905 101.455 113.905 101.625 ;
        RECT 114.195 101.455 116.195 101.625 ;
        RECT 116.485 101.455 118.485 101.625 ;
        RECT 118.775 101.455 120.775 101.625 ;
        RECT 121.065 101.455 123.065 101.625 ;
        RECT 123.355 101.455 125.355 101.625 ;
        RECT 125.645 101.455 127.645 101.625 ;
        RECT 109.385 93.200 109.555 101.240 ;
        RECT 111.675 93.200 111.845 101.240 ;
        RECT 113.965 93.200 114.135 101.240 ;
        RECT 116.255 93.200 116.425 101.240 ;
        RECT 118.545 93.200 118.715 101.240 ;
        RECT 120.835 93.200 121.005 101.240 ;
        RECT 123.125 93.200 123.295 101.240 ;
        RECT 125.415 93.200 125.585 101.240 ;
        RECT 127.705 93.200 127.875 101.240 ;
        RECT 109.615 92.815 111.615 92.985 ;
        RECT 111.905 92.815 113.905 92.985 ;
        RECT 114.195 92.815 116.195 92.985 ;
        RECT 116.485 92.815 118.485 92.985 ;
        RECT 118.775 92.815 120.775 92.985 ;
        RECT 121.065 92.815 123.065 92.985 ;
        RECT 123.355 92.815 125.355 92.985 ;
        RECT 125.645 92.815 127.645 92.985 ;
        RECT 128.375 92.295 128.905 102.145 ;
        RECT 10.055 92.125 128.905 92.295 ;
        RECT 10.055 82.275 10.585 92.125 ;
        RECT 11.315 91.435 13.315 91.605 ;
        RECT 13.605 91.435 15.605 91.605 ;
        RECT 15.895 91.435 17.895 91.605 ;
        RECT 18.185 91.435 20.185 91.605 ;
        RECT 20.475 91.435 22.475 91.605 ;
        RECT 22.765 91.435 24.765 91.605 ;
        RECT 25.055 91.435 27.055 91.605 ;
        RECT 27.345 91.435 29.345 91.605 ;
        RECT 11.085 83.180 11.255 91.220 ;
        RECT 13.375 83.180 13.545 91.220 ;
        RECT 15.665 83.180 15.835 91.220 ;
        RECT 17.955 83.180 18.125 91.220 ;
        RECT 20.245 83.180 20.415 91.220 ;
        RECT 22.535 83.180 22.705 91.220 ;
        RECT 24.825 83.180 24.995 91.220 ;
        RECT 27.115 83.180 27.285 91.220 ;
        RECT 29.405 83.180 29.575 91.220 ;
        RECT 11.315 82.795 13.315 82.965 ;
        RECT 13.605 82.795 15.605 82.965 ;
        RECT 15.895 82.795 17.895 82.965 ;
        RECT 18.185 82.795 20.185 82.965 ;
        RECT 20.475 82.795 22.475 82.965 ;
        RECT 22.765 82.795 24.765 82.965 ;
        RECT 25.055 82.795 27.055 82.965 ;
        RECT 27.345 82.795 29.345 82.965 ;
        RECT 30.075 82.275 30.245 92.125 ;
        RECT 30.975 91.435 32.975 91.605 ;
        RECT 33.265 91.435 35.265 91.605 ;
        RECT 35.555 91.435 37.555 91.605 ;
        RECT 37.845 91.435 39.845 91.605 ;
        RECT 40.135 91.435 42.135 91.605 ;
        RECT 42.425 91.435 44.425 91.605 ;
        RECT 44.715 91.435 46.715 91.605 ;
        RECT 47.005 91.435 49.005 91.605 ;
        RECT 30.745 83.180 30.915 91.220 ;
        RECT 33.035 83.180 33.205 91.220 ;
        RECT 35.325 83.180 35.495 91.220 ;
        RECT 37.615 83.180 37.785 91.220 ;
        RECT 39.905 83.180 40.075 91.220 ;
        RECT 42.195 83.180 42.365 91.220 ;
        RECT 44.485 83.180 44.655 91.220 ;
        RECT 46.775 83.180 46.945 91.220 ;
        RECT 49.065 83.180 49.235 91.220 ;
        RECT 30.975 82.795 32.975 82.965 ;
        RECT 33.265 82.795 35.265 82.965 ;
        RECT 35.555 82.795 37.555 82.965 ;
        RECT 37.845 82.795 39.845 82.965 ;
        RECT 40.135 82.795 42.135 82.965 ;
        RECT 42.425 82.795 44.425 82.965 ;
        RECT 44.715 82.795 46.715 82.965 ;
        RECT 47.005 82.795 49.005 82.965 ;
        RECT 49.735 82.275 49.905 92.125 ;
        RECT 50.635 91.435 52.635 91.605 ;
        RECT 52.925 91.435 54.925 91.605 ;
        RECT 55.215 91.435 57.215 91.605 ;
        RECT 57.505 91.435 59.505 91.605 ;
        RECT 59.795 91.435 61.795 91.605 ;
        RECT 62.085 91.435 64.085 91.605 ;
        RECT 64.375 91.435 66.375 91.605 ;
        RECT 66.665 91.435 68.665 91.605 ;
        RECT 50.405 83.180 50.575 91.220 ;
        RECT 52.695 83.180 52.865 91.220 ;
        RECT 54.985 83.180 55.155 91.220 ;
        RECT 57.275 83.180 57.445 91.220 ;
        RECT 59.565 83.180 59.735 91.220 ;
        RECT 61.855 83.180 62.025 91.220 ;
        RECT 64.145 83.180 64.315 91.220 ;
        RECT 66.435 83.180 66.605 91.220 ;
        RECT 68.725 83.180 68.895 91.220 ;
        RECT 50.635 82.795 52.635 82.965 ;
        RECT 52.925 82.795 54.925 82.965 ;
        RECT 55.215 82.795 57.215 82.965 ;
        RECT 57.505 82.795 59.505 82.965 ;
        RECT 59.795 82.795 61.795 82.965 ;
        RECT 62.085 82.795 64.085 82.965 ;
        RECT 64.375 82.795 66.375 82.965 ;
        RECT 66.665 82.795 68.665 82.965 ;
        RECT 69.395 82.275 69.565 92.125 ;
        RECT 70.295 91.435 72.295 91.605 ;
        RECT 72.585 91.435 74.585 91.605 ;
        RECT 74.875 91.435 76.875 91.605 ;
        RECT 77.165 91.435 79.165 91.605 ;
        RECT 79.455 91.435 81.455 91.605 ;
        RECT 81.745 91.435 83.745 91.605 ;
        RECT 84.035 91.435 86.035 91.605 ;
        RECT 86.325 91.435 88.325 91.605 ;
        RECT 70.065 83.180 70.235 91.220 ;
        RECT 72.355 83.180 72.525 91.220 ;
        RECT 74.645 83.180 74.815 91.220 ;
        RECT 76.935 83.180 77.105 91.220 ;
        RECT 79.225 83.180 79.395 91.220 ;
        RECT 81.515 83.180 81.685 91.220 ;
        RECT 83.805 83.180 83.975 91.220 ;
        RECT 86.095 83.180 86.265 91.220 ;
        RECT 88.385 83.180 88.555 91.220 ;
        RECT 70.295 82.795 72.295 82.965 ;
        RECT 72.585 82.795 74.585 82.965 ;
        RECT 74.875 82.795 76.875 82.965 ;
        RECT 77.165 82.795 79.165 82.965 ;
        RECT 79.455 82.795 81.455 82.965 ;
        RECT 81.745 82.795 83.745 82.965 ;
        RECT 84.035 82.795 86.035 82.965 ;
        RECT 86.325 82.795 88.325 82.965 ;
        RECT 89.055 82.275 89.225 92.125 ;
        RECT 89.955 91.435 91.955 91.605 ;
        RECT 92.245 91.435 94.245 91.605 ;
        RECT 94.535 91.435 96.535 91.605 ;
        RECT 96.825 91.435 98.825 91.605 ;
        RECT 99.115 91.435 101.115 91.605 ;
        RECT 101.405 91.435 103.405 91.605 ;
        RECT 103.695 91.435 105.695 91.605 ;
        RECT 105.985 91.435 107.985 91.605 ;
        RECT 89.725 83.180 89.895 91.220 ;
        RECT 92.015 83.180 92.185 91.220 ;
        RECT 94.305 83.180 94.475 91.220 ;
        RECT 96.595 83.180 96.765 91.220 ;
        RECT 98.885 83.180 99.055 91.220 ;
        RECT 101.175 83.180 101.345 91.220 ;
        RECT 103.465 83.180 103.635 91.220 ;
        RECT 105.755 83.180 105.925 91.220 ;
        RECT 108.045 83.180 108.215 91.220 ;
        RECT 89.955 82.795 91.955 82.965 ;
        RECT 92.245 82.795 94.245 82.965 ;
        RECT 94.535 82.795 96.535 82.965 ;
        RECT 96.825 82.795 98.825 82.965 ;
        RECT 99.115 82.795 101.115 82.965 ;
        RECT 101.405 82.795 103.405 82.965 ;
        RECT 103.695 82.795 105.695 82.965 ;
        RECT 105.985 82.795 107.985 82.965 ;
        RECT 108.715 82.275 108.885 92.125 ;
        RECT 109.615 91.435 111.615 91.605 ;
        RECT 111.905 91.435 113.905 91.605 ;
        RECT 114.195 91.435 116.195 91.605 ;
        RECT 116.485 91.435 118.485 91.605 ;
        RECT 118.775 91.435 120.775 91.605 ;
        RECT 121.065 91.435 123.065 91.605 ;
        RECT 123.355 91.435 125.355 91.605 ;
        RECT 125.645 91.435 127.645 91.605 ;
        RECT 109.385 83.180 109.555 91.220 ;
        RECT 111.675 83.180 111.845 91.220 ;
        RECT 113.965 83.180 114.135 91.220 ;
        RECT 116.255 83.180 116.425 91.220 ;
        RECT 118.545 83.180 118.715 91.220 ;
        RECT 120.835 83.180 121.005 91.220 ;
        RECT 123.125 83.180 123.295 91.220 ;
        RECT 125.415 83.180 125.585 91.220 ;
        RECT 127.705 83.180 127.875 91.220 ;
        RECT 109.615 82.795 111.615 82.965 ;
        RECT 111.905 82.795 113.905 82.965 ;
        RECT 114.195 82.795 116.195 82.965 ;
        RECT 116.485 82.795 118.485 82.965 ;
        RECT 118.775 82.795 120.775 82.965 ;
        RECT 121.065 82.795 123.065 82.965 ;
        RECT 123.355 82.795 125.355 82.965 ;
        RECT 125.645 82.795 127.645 82.965 ;
        RECT 128.375 82.275 128.905 92.125 ;
        RECT 10.055 82.105 128.905 82.275 ;
        RECT 10.055 72.255 10.585 82.105 ;
        RECT 11.315 81.415 13.315 81.585 ;
        RECT 13.605 81.415 15.605 81.585 ;
        RECT 15.895 81.415 17.895 81.585 ;
        RECT 18.185 81.415 20.185 81.585 ;
        RECT 20.475 81.415 22.475 81.585 ;
        RECT 22.765 81.415 24.765 81.585 ;
        RECT 25.055 81.415 27.055 81.585 ;
        RECT 27.345 81.415 29.345 81.585 ;
        RECT 11.085 73.160 11.255 81.200 ;
        RECT 13.375 73.160 13.545 81.200 ;
        RECT 15.665 73.160 15.835 81.200 ;
        RECT 17.955 73.160 18.125 81.200 ;
        RECT 20.245 73.160 20.415 81.200 ;
        RECT 22.535 73.160 22.705 81.200 ;
        RECT 24.825 73.160 24.995 81.200 ;
        RECT 27.115 73.160 27.285 81.200 ;
        RECT 29.405 73.160 29.575 81.200 ;
        RECT 11.315 72.775 13.315 72.945 ;
        RECT 13.605 72.775 15.605 72.945 ;
        RECT 15.895 72.775 17.895 72.945 ;
        RECT 18.185 72.775 20.185 72.945 ;
        RECT 20.475 72.775 22.475 72.945 ;
        RECT 22.765 72.775 24.765 72.945 ;
        RECT 25.055 72.775 27.055 72.945 ;
        RECT 27.345 72.775 29.345 72.945 ;
        RECT 30.075 72.255 30.245 82.105 ;
        RECT 30.975 81.415 32.975 81.585 ;
        RECT 33.265 81.415 35.265 81.585 ;
        RECT 35.555 81.415 37.555 81.585 ;
        RECT 37.845 81.415 39.845 81.585 ;
        RECT 40.135 81.415 42.135 81.585 ;
        RECT 42.425 81.415 44.425 81.585 ;
        RECT 44.715 81.415 46.715 81.585 ;
        RECT 47.005 81.415 49.005 81.585 ;
        RECT 30.745 73.160 30.915 81.200 ;
        RECT 33.035 73.160 33.205 81.200 ;
        RECT 35.325 73.160 35.495 81.200 ;
        RECT 37.615 73.160 37.785 81.200 ;
        RECT 39.905 73.160 40.075 81.200 ;
        RECT 42.195 73.160 42.365 81.200 ;
        RECT 44.485 73.160 44.655 81.200 ;
        RECT 46.775 73.160 46.945 81.200 ;
        RECT 49.065 73.160 49.235 81.200 ;
        RECT 30.975 72.775 32.975 72.945 ;
        RECT 33.265 72.775 35.265 72.945 ;
        RECT 35.555 72.775 37.555 72.945 ;
        RECT 37.845 72.775 39.845 72.945 ;
        RECT 40.135 72.775 42.135 72.945 ;
        RECT 42.425 72.775 44.425 72.945 ;
        RECT 44.715 72.775 46.715 72.945 ;
        RECT 47.005 72.775 49.005 72.945 ;
        RECT 49.735 72.255 49.905 82.105 ;
        RECT 50.635 81.415 52.635 81.585 ;
        RECT 52.925 81.415 54.925 81.585 ;
        RECT 55.215 81.415 57.215 81.585 ;
        RECT 57.505 81.415 59.505 81.585 ;
        RECT 59.795 81.415 61.795 81.585 ;
        RECT 62.085 81.415 64.085 81.585 ;
        RECT 64.375 81.415 66.375 81.585 ;
        RECT 66.665 81.415 68.665 81.585 ;
        RECT 50.405 73.160 50.575 81.200 ;
        RECT 52.695 73.160 52.865 81.200 ;
        RECT 54.985 73.160 55.155 81.200 ;
        RECT 57.275 73.160 57.445 81.200 ;
        RECT 59.565 73.160 59.735 81.200 ;
        RECT 61.855 73.160 62.025 81.200 ;
        RECT 64.145 73.160 64.315 81.200 ;
        RECT 66.435 73.160 66.605 81.200 ;
        RECT 68.725 73.160 68.895 81.200 ;
        RECT 50.635 72.775 52.635 72.945 ;
        RECT 52.925 72.775 54.925 72.945 ;
        RECT 55.215 72.775 57.215 72.945 ;
        RECT 57.505 72.775 59.505 72.945 ;
        RECT 59.795 72.775 61.795 72.945 ;
        RECT 62.085 72.775 64.085 72.945 ;
        RECT 64.375 72.775 66.375 72.945 ;
        RECT 66.665 72.775 68.665 72.945 ;
        RECT 69.395 72.255 69.565 82.105 ;
        RECT 70.295 81.415 72.295 81.585 ;
        RECT 72.585 81.415 74.585 81.585 ;
        RECT 74.875 81.415 76.875 81.585 ;
        RECT 77.165 81.415 79.165 81.585 ;
        RECT 79.455 81.415 81.455 81.585 ;
        RECT 81.745 81.415 83.745 81.585 ;
        RECT 84.035 81.415 86.035 81.585 ;
        RECT 86.325 81.415 88.325 81.585 ;
        RECT 70.065 73.160 70.235 81.200 ;
        RECT 72.355 73.160 72.525 81.200 ;
        RECT 74.645 73.160 74.815 81.200 ;
        RECT 76.935 73.160 77.105 81.200 ;
        RECT 79.225 73.160 79.395 81.200 ;
        RECT 81.515 73.160 81.685 81.200 ;
        RECT 83.805 73.160 83.975 81.200 ;
        RECT 86.095 73.160 86.265 81.200 ;
        RECT 88.385 73.160 88.555 81.200 ;
        RECT 70.295 72.775 72.295 72.945 ;
        RECT 72.585 72.775 74.585 72.945 ;
        RECT 74.875 72.775 76.875 72.945 ;
        RECT 77.165 72.775 79.165 72.945 ;
        RECT 79.455 72.775 81.455 72.945 ;
        RECT 81.745 72.775 83.745 72.945 ;
        RECT 84.035 72.775 86.035 72.945 ;
        RECT 86.325 72.775 88.325 72.945 ;
        RECT 89.055 72.255 89.225 82.105 ;
        RECT 89.955 81.415 91.955 81.585 ;
        RECT 92.245 81.415 94.245 81.585 ;
        RECT 94.535 81.415 96.535 81.585 ;
        RECT 96.825 81.415 98.825 81.585 ;
        RECT 99.115 81.415 101.115 81.585 ;
        RECT 101.405 81.415 103.405 81.585 ;
        RECT 103.695 81.415 105.695 81.585 ;
        RECT 105.985 81.415 107.985 81.585 ;
        RECT 89.725 73.160 89.895 81.200 ;
        RECT 92.015 73.160 92.185 81.200 ;
        RECT 94.305 73.160 94.475 81.200 ;
        RECT 96.595 73.160 96.765 81.200 ;
        RECT 98.885 73.160 99.055 81.200 ;
        RECT 101.175 73.160 101.345 81.200 ;
        RECT 103.465 73.160 103.635 81.200 ;
        RECT 105.755 73.160 105.925 81.200 ;
        RECT 108.045 73.160 108.215 81.200 ;
        RECT 89.955 72.775 91.955 72.945 ;
        RECT 92.245 72.775 94.245 72.945 ;
        RECT 94.535 72.775 96.535 72.945 ;
        RECT 96.825 72.775 98.825 72.945 ;
        RECT 99.115 72.775 101.115 72.945 ;
        RECT 101.405 72.775 103.405 72.945 ;
        RECT 103.695 72.775 105.695 72.945 ;
        RECT 105.985 72.775 107.985 72.945 ;
        RECT 108.715 72.255 108.885 82.105 ;
        RECT 109.615 81.415 111.615 81.585 ;
        RECT 111.905 81.415 113.905 81.585 ;
        RECT 114.195 81.415 116.195 81.585 ;
        RECT 116.485 81.415 118.485 81.585 ;
        RECT 118.775 81.415 120.775 81.585 ;
        RECT 121.065 81.415 123.065 81.585 ;
        RECT 123.355 81.415 125.355 81.585 ;
        RECT 125.645 81.415 127.645 81.585 ;
        RECT 109.385 73.160 109.555 81.200 ;
        RECT 111.675 73.160 111.845 81.200 ;
        RECT 113.965 73.160 114.135 81.200 ;
        RECT 116.255 73.160 116.425 81.200 ;
        RECT 118.545 73.160 118.715 81.200 ;
        RECT 120.835 73.160 121.005 81.200 ;
        RECT 123.125 73.160 123.295 81.200 ;
        RECT 125.415 73.160 125.585 81.200 ;
        RECT 127.705 73.160 127.875 81.200 ;
        RECT 109.615 72.775 111.615 72.945 ;
        RECT 111.905 72.775 113.905 72.945 ;
        RECT 114.195 72.775 116.195 72.945 ;
        RECT 116.485 72.775 118.485 72.945 ;
        RECT 118.775 72.775 120.775 72.945 ;
        RECT 121.065 72.775 123.065 72.945 ;
        RECT 123.355 72.775 125.355 72.945 ;
        RECT 125.645 72.775 127.645 72.945 ;
        RECT 128.375 72.255 128.905 82.105 ;
        RECT 10.055 72.085 128.905 72.255 ;
        RECT 10.055 62.235 10.585 72.085 ;
        RECT 11.315 71.395 13.315 71.565 ;
        RECT 13.605 71.395 15.605 71.565 ;
        RECT 15.895 71.395 17.895 71.565 ;
        RECT 18.185 71.395 20.185 71.565 ;
        RECT 20.475 71.395 22.475 71.565 ;
        RECT 22.765 71.395 24.765 71.565 ;
        RECT 25.055 71.395 27.055 71.565 ;
        RECT 27.345 71.395 29.345 71.565 ;
        RECT 11.085 63.140 11.255 71.180 ;
        RECT 13.375 63.140 13.545 71.180 ;
        RECT 15.665 63.140 15.835 71.180 ;
        RECT 17.955 63.140 18.125 71.180 ;
        RECT 20.245 63.140 20.415 71.180 ;
        RECT 22.535 63.140 22.705 71.180 ;
        RECT 24.825 63.140 24.995 71.180 ;
        RECT 27.115 63.140 27.285 71.180 ;
        RECT 29.405 63.140 29.575 71.180 ;
        RECT 11.315 62.755 13.315 62.925 ;
        RECT 13.605 62.755 15.605 62.925 ;
        RECT 15.895 62.755 17.895 62.925 ;
        RECT 18.185 62.755 20.185 62.925 ;
        RECT 20.475 62.755 22.475 62.925 ;
        RECT 22.765 62.755 24.765 62.925 ;
        RECT 25.055 62.755 27.055 62.925 ;
        RECT 27.345 62.755 29.345 62.925 ;
        RECT 30.075 62.235 30.245 72.085 ;
        RECT 30.975 71.395 32.975 71.565 ;
        RECT 33.265 71.395 35.265 71.565 ;
        RECT 35.555 71.395 37.555 71.565 ;
        RECT 37.845 71.395 39.845 71.565 ;
        RECT 40.135 71.395 42.135 71.565 ;
        RECT 42.425 71.395 44.425 71.565 ;
        RECT 44.715 71.395 46.715 71.565 ;
        RECT 47.005 71.395 49.005 71.565 ;
        RECT 30.745 63.140 30.915 71.180 ;
        RECT 33.035 63.140 33.205 71.180 ;
        RECT 35.325 63.140 35.495 71.180 ;
        RECT 37.615 63.140 37.785 71.180 ;
        RECT 39.905 63.140 40.075 71.180 ;
        RECT 42.195 63.140 42.365 71.180 ;
        RECT 44.485 63.140 44.655 71.180 ;
        RECT 46.775 63.140 46.945 71.180 ;
        RECT 49.065 63.140 49.235 71.180 ;
        RECT 30.975 62.755 32.975 62.925 ;
        RECT 33.265 62.755 35.265 62.925 ;
        RECT 35.555 62.755 37.555 62.925 ;
        RECT 37.845 62.755 39.845 62.925 ;
        RECT 40.135 62.755 42.135 62.925 ;
        RECT 42.425 62.755 44.425 62.925 ;
        RECT 44.715 62.755 46.715 62.925 ;
        RECT 47.005 62.755 49.005 62.925 ;
        RECT 49.735 62.235 49.905 72.085 ;
        RECT 50.635 71.395 52.635 71.565 ;
        RECT 52.925 71.395 54.925 71.565 ;
        RECT 55.215 71.395 57.215 71.565 ;
        RECT 57.505 71.395 59.505 71.565 ;
        RECT 59.795 71.395 61.795 71.565 ;
        RECT 62.085 71.395 64.085 71.565 ;
        RECT 64.375 71.395 66.375 71.565 ;
        RECT 66.665 71.395 68.665 71.565 ;
        RECT 50.405 63.140 50.575 71.180 ;
        RECT 52.695 63.140 52.865 71.180 ;
        RECT 54.985 63.140 55.155 71.180 ;
        RECT 57.275 63.140 57.445 71.180 ;
        RECT 59.565 63.140 59.735 71.180 ;
        RECT 61.855 63.140 62.025 71.180 ;
        RECT 64.145 63.140 64.315 71.180 ;
        RECT 66.435 63.140 66.605 71.180 ;
        RECT 68.725 63.140 68.895 71.180 ;
        RECT 50.635 62.755 52.635 62.925 ;
        RECT 52.925 62.755 54.925 62.925 ;
        RECT 55.215 62.755 57.215 62.925 ;
        RECT 57.505 62.755 59.505 62.925 ;
        RECT 59.795 62.755 61.795 62.925 ;
        RECT 62.085 62.755 64.085 62.925 ;
        RECT 64.375 62.755 66.375 62.925 ;
        RECT 66.665 62.755 68.665 62.925 ;
        RECT 69.395 62.235 69.565 72.085 ;
        RECT 70.295 71.395 72.295 71.565 ;
        RECT 72.585 71.395 74.585 71.565 ;
        RECT 74.875 71.395 76.875 71.565 ;
        RECT 77.165 71.395 79.165 71.565 ;
        RECT 79.455 71.395 81.455 71.565 ;
        RECT 81.745 71.395 83.745 71.565 ;
        RECT 84.035 71.395 86.035 71.565 ;
        RECT 86.325 71.395 88.325 71.565 ;
        RECT 70.065 63.140 70.235 71.180 ;
        RECT 72.355 63.140 72.525 71.180 ;
        RECT 74.645 63.140 74.815 71.180 ;
        RECT 76.935 63.140 77.105 71.180 ;
        RECT 79.225 63.140 79.395 71.180 ;
        RECT 81.515 63.140 81.685 71.180 ;
        RECT 83.805 63.140 83.975 71.180 ;
        RECT 86.095 63.140 86.265 71.180 ;
        RECT 88.385 63.140 88.555 71.180 ;
        RECT 70.295 62.755 72.295 62.925 ;
        RECT 72.585 62.755 74.585 62.925 ;
        RECT 74.875 62.755 76.875 62.925 ;
        RECT 77.165 62.755 79.165 62.925 ;
        RECT 79.455 62.755 81.455 62.925 ;
        RECT 81.745 62.755 83.745 62.925 ;
        RECT 84.035 62.755 86.035 62.925 ;
        RECT 86.325 62.755 88.325 62.925 ;
        RECT 89.055 62.235 89.225 72.085 ;
        RECT 89.955 71.395 91.955 71.565 ;
        RECT 92.245 71.395 94.245 71.565 ;
        RECT 94.535 71.395 96.535 71.565 ;
        RECT 96.825 71.395 98.825 71.565 ;
        RECT 99.115 71.395 101.115 71.565 ;
        RECT 101.405 71.395 103.405 71.565 ;
        RECT 103.695 71.395 105.695 71.565 ;
        RECT 105.985 71.395 107.985 71.565 ;
        RECT 89.725 63.140 89.895 71.180 ;
        RECT 92.015 63.140 92.185 71.180 ;
        RECT 94.305 63.140 94.475 71.180 ;
        RECT 96.595 63.140 96.765 71.180 ;
        RECT 98.885 63.140 99.055 71.180 ;
        RECT 101.175 63.140 101.345 71.180 ;
        RECT 103.465 63.140 103.635 71.180 ;
        RECT 105.755 63.140 105.925 71.180 ;
        RECT 108.045 63.140 108.215 71.180 ;
        RECT 89.955 62.755 91.955 62.925 ;
        RECT 92.245 62.755 94.245 62.925 ;
        RECT 94.535 62.755 96.535 62.925 ;
        RECT 96.825 62.755 98.825 62.925 ;
        RECT 99.115 62.755 101.115 62.925 ;
        RECT 101.405 62.755 103.405 62.925 ;
        RECT 103.695 62.755 105.695 62.925 ;
        RECT 105.985 62.755 107.985 62.925 ;
        RECT 108.715 62.235 108.885 72.085 ;
        RECT 109.615 71.395 111.615 71.565 ;
        RECT 111.905 71.395 113.905 71.565 ;
        RECT 114.195 71.395 116.195 71.565 ;
        RECT 116.485 71.395 118.485 71.565 ;
        RECT 118.775 71.395 120.775 71.565 ;
        RECT 121.065 71.395 123.065 71.565 ;
        RECT 123.355 71.395 125.355 71.565 ;
        RECT 125.645 71.395 127.645 71.565 ;
        RECT 109.385 63.140 109.555 71.180 ;
        RECT 111.675 63.140 111.845 71.180 ;
        RECT 113.965 63.140 114.135 71.180 ;
        RECT 116.255 63.140 116.425 71.180 ;
        RECT 118.545 63.140 118.715 71.180 ;
        RECT 120.835 63.140 121.005 71.180 ;
        RECT 123.125 63.140 123.295 71.180 ;
        RECT 125.415 63.140 125.585 71.180 ;
        RECT 127.705 63.140 127.875 71.180 ;
        RECT 109.615 62.755 111.615 62.925 ;
        RECT 111.905 62.755 113.905 62.925 ;
        RECT 114.195 62.755 116.195 62.925 ;
        RECT 116.485 62.755 118.485 62.925 ;
        RECT 118.775 62.755 120.775 62.925 ;
        RECT 121.065 62.755 123.065 62.925 ;
        RECT 123.355 62.755 125.355 62.925 ;
        RECT 125.645 62.755 127.645 62.925 ;
        RECT 128.375 62.235 128.905 72.085 ;
        RECT 10.055 62.065 128.905 62.235 ;
        RECT 10.055 52.215 10.585 62.065 ;
        RECT 11.315 61.375 13.315 61.545 ;
        RECT 13.605 61.375 15.605 61.545 ;
        RECT 15.895 61.375 17.895 61.545 ;
        RECT 18.185 61.375 20.185 61.545 ;
        RECT 20.475 61.375 22.475 61.545 ;
        RECT 22.765 61.375 24.765 61.545 ;
        RECT 25.055 61.375 27.055 61.545 ;
        RECT 27.345 61.375 29.345 61.545 ;
        RECT 11.085 53.120 11.255 61.160 ;
        RECT 13.375 53.120 13.545 61.160 ;
        RECT 15.665 53.120 15.835 61.160 ;
        RECT 17.955 53.120 18.125 61.160 ;
        RECT 20.245 53.120 20.415 61.160 ;
        RECT 22.535 53.120 22.705 61.160 ;
        RECT 24.825 53.120 24.995 61.160 ;
        RECT 27.115 53.120 27.285 61.160 ;
        RECT 29.405 53.120 29.575 61.160 ;
        RECT 11.315 52.735 13.315 52.905 ;
        RECT 13.605 52.735 15.605 52.905 ;
        RECT 15.895 52.735 17.895 52.905 ;
        RECT 18.185 52.735 20.185 52.905 ;
        RECT 20.475 52.735 22.475 52.905 ;
        RECT 22.765 52.735 24.765 52.905 ;
        RECT 25.055 52.735 27.055 52.905 ;
        RECT 27.345 52.735 29.345 52.905 ;
        RECT 30.075 52.215 30.245 62.065 ;
        RECT 30.975 61.375 32.975 61.545 ;
        RECT 33.265 61.375 35.265 61.545 ;
        RECT 35.555 61.375 37.555 61.545 ;
        RECT 37.845 61.375 39.845 61.545 ;
        RECT 40.135 61.375 42.135 61.545 ;
        RECT 42.425 61.375 44.425 61.545 ;
        RECT 44.715 61.375 46.715 61.545 ;
        RECT 47.005 61.375 49.005 61.545 ;
        RECT 30.745 53.120 30.915 61.160 ;
        RECT 33.035 53.120 33.205 61.160 ;
        RECT 35.325 53.120 35.495 61.160 ;
        RECT 37.615 53.120 37.785 61.160 ;
        RECT 39.905 53.120 40.075 61.160 ;
        RECT 42.195 53.120 42.365 61.160 ;
        RECT 44.485 53.120 44.655 61.160 ;
        RECT 46.775 53.120 46.945 61.160 ;
        RECT 49.065 53.120 49.235 61.160 ;
        RECT 30.975 52.735 32.975 52.905 ;
        RECT 33.265 52.735 35.265 52.905 ;
        RECT 35.555 52.735 37.555 52.905 ;
        RECT 37.845 52.735 39.845 52.905 ;
        RECT 40.135 52.735 42.135 52.905 ;
        RECT 42.425 52.735 44.425 52.905 ;
        RECT 44.715 52.735 46.715 52.905 ;
        RECT 47.005 52.735 49.005 52.905 ;
        RECT 49.735 52.215 49.905 62.065 ;
        RECT 50.635 61.375 52.635 61.545 ;
        RECT 52.925 61.375 54.925 61.545 ;
        RECT 55.215 61.375 57.215 61.545 ;
        RECT 57.505 61.375 59.505 61.545 ;
        RECT 59.795 61.375 61.795 61.545 ;
        RECT 62.085 61.375 64.085 61.545 ;
        RECT 64.375 61.375 66.375 61.545 ;
        RECT 66.665 61.375 68.665 61.545 ;
        RECT 50.405 53.120 50.575 61.160 ;
        RECT 52.695 53.120 52.865 61.160 ;
        RECT 54.985 53.120 55.155 61.160 ;
        RECT 57.275 53.120 57.445 61.160 ;
        RECT 59.565 53.120 59.735 61.160 ;
        RECT 61.855 53.120 62.025 61.160 ;
        RECT 64.145 53.120 64.315 61.160 ;
        RECT 66.435 53.120 66.605 61.160 ;
        RECT 68.725 53.120 68.895 61.160 ;
        RECT 50.635 52.735 52.635 52.905 ;
        RECT 52.925 52.735 54.925 52.905 ;
        RECT 55.215 52.735 57.215 52.905 ;
        RECT 57.505 52.735 59.505 52.905 ;
        RECT 59.795 52.735 61.795 52.905 ;
        RECT 62.085 52.735 64.085 52.905 ;
        RECT 64.375 52.735 66.375 52.905 ;
        RECT 66.665 52.735 68.665 52.905 ;
        RECT 69.395 52.215 69.565 62.065 ;
        RECT 70.295 61.375 72.295 61.545 ;
        RECT 72.585 61.375 74.585 61.545 ;
        RECT 74.875 61.375 76.875 61.545 ;
        RECT 77.165 61.375 79.165 61.545 ;
        RECT 79.455 61.375 81.455 61.545 ;
        RECT 81.745 61.375 83.745 61.545 ;
        RECT 84.035 61.375 86.035 61.545 ;
        RECT 86.325 61.375 88.325 61.545 ;
        RECT 70.065 53.120 70.235 61.160 ;
        RECT 72.355 53.120 72.525 61.160 ;
        RECT 74.645 53.120 74.815 61.160 ;
        RECT 76.935 53.120 77.105 61.160 ;
        RECT 79.225 53.120 79.395 61.160 ;
        RECT 81.515 53.120 81.685 61.160 ;
        RECT 83.805 53.120 83.975 61.160 ;
        RECT 86.095 53.120 86.265 61.160 ;
        RECT 88.385 53.120 88.555 61.160 ;
        RECT 70.295 52.735 72.295 52.905 ;
        RECT 72.585 52.735 74.585 52.905 ;
        RECT 74.875 52.735 76.875 52.905 ;
        RECT 77.165 52.735 79.165 52.905 ;
        RECT 79.455 52.735 81.455 52.905 ;
        RECT 81.745 52.735 83.745 52.905 ;
        RECT 84.035 52.735 86.035 52.905 ;
        RECT 86.325 52.735 88.325 52.905 ;
        RECT 89.055 52.215 89.225 62.065 ;
        RECT 89.955 61.375 91.955 61.545 ;
        RECT 92.245 61.375 94.245 61.545 ;
        RECT 94.535 61.375 96.535 61.545 ;
        RECT 96.825 61.375 98.825 61.545 ;
        RECT 99.115 61.375 101.115 61.545 ;
        RECT 101.405 61.375 103.405 61.545 ;
        RECT 103.695 61.375 105.695 61.545 ;
        RECT 105.985 61.375 107.985 61.545 ;
        RECT 89.725 53.120 89.895 61.160 ;
        RECT 92.015 53.120 92.185 61.160 ;
        RECT 94.305 53.120 94.475 61.160 ;
        RECT 96.595 53.120 96.765 61.160 ;
        RECT 98.885 53.120 99.055 61.160 ;
        RECT 101.175 53.120 101.345 61.160 ;
        RECT 103.465 53.120 103.635 61.160 ;
        RECT 105.755 53.120 105.925 61.160 ;
        RECT 108.045 53.120 108.215 61.160 ;
        RECT 89.955 52.735 91.955 52.905 ;
        RECT 92.245 52.735 94.245 52.905 ;
        RECT 94.535 52.735 96.535 52.905 ;
        RECT 96.825 52.735 98.825 52.905 ;
        RECT 99.115 52.735 101.115 52.905 ;
        RECT 101.405 52.735 103.405 52.905 ;
        RECT 103.695 52.735 105.695 52.905 ;
        RECT 105.985 52.735 107.985 52.905 ;
        RECT 108.715 52.215 108.885 62.065 ;
        RECT 109.615 61.375 111.615 61.545 ;
        RECT 111.905 61.375 113.905 61.545 ;
        RECT 114.195 61.375 116.195 61.545 ;
        RECT 116.485 61.375 118.485 61.545 ;
        RECT 118.775 61.375 120.775 61.545 ;
        RECT 121.065 61.375 123.065 61.545 ;
        RECT 123.355 61.375 125.355 61.545 ;
        RECT 125.645 61.375 127.645 61.545 ;
        RECT 109.385 53.120 109.555 61.160 ;
        RECT 111.675 53.120 111.845 61.160 ;
        RECT 113.965 53.120 114.135 61.160 ;
        RECT 116.255 53.120 116.425 61.160 ;
        RECT 118.545 53.120 118.715 61.160 ;
        RECT 120.835 53.120 121.005 61.160 ;
        RECT 123.125 53.120 123.295 61.160 ;
        RECT 125.415 53.120 125.585 61.160 ;
        RECT 127.705 53.120 127.875 61.160 ;
        RECT 109.615 52.735 111.615 52.905 ;
        RECT 111.905 52.735 113.905 52.905 ;
        RECT 114.195 52.735 116.195 52.905 ;
        RECT 116.485 52.735 118.485 52.905 ;
        RECT 118.775 52.735 120.775 52.905 ;
        RECT 121.065 52.735 123.065 52.905 ;
        RECT 123.355 52.735 125.355 52.905 ;
        RECT 125.645 52.735 127.645 52.905 ;
        RECT 128.375 52.215 128.905 62.065 ;
        RECT 10.055 52.045 128.905 52.215 ;
        RECT 10.055 42.195 10.585 52.045 ;
        RECT 11.315 51.355 13.315 51.525 ;
        RECT 13.605 51.355 15.605 51.525 ;
        RECT 15.895 51.355 17.895 51.525 ;
        RECT 18.185 51.355 20.185 51.525 ;
        RECT 20.475 51.355 22.475 51.525 ;
        RECT 22.765 51.355 24.765 51.525 ;
        RECT 25.055 51.355 27.055 51.525 ;
        RECT 27.345 51.355 29.345 51.525 ;
        RECT 11.085 43.100 11.255 51.140 ;
        RECT 13.375 43.100 13.545 51.140 ;
        RECT 15.665 43.100 15.835 51.140 ;
        RECT 17.955 43.100 18.125 51.140 ;
        RECT 20.245 43.100 20.415 51.140 ;
        RECT 22.535 43.100 22.705 51.140 ;
        RECT 24.825 43.100 24.995 51.140 ;
        RECT 27.115 43.100 27.285 51.140 ;
        RECT 29.405 43.100 29.575 51.140 ;
        RECT 11.315 42.715 13.315 42.885 ;
        RECT 13.605 42.715 15.605 42.885 ;
        RECT 15.895 42.715 17.895 42.885 ;
        RECT 18.185 42.715 20.185 42.885 ;
        RECT 20.475 42.715 22.475 42.885 ;
        RECT 22.765 42.715 24.765 42.885 ;
        RECT 25.055 42.715 27.055 42.885 ;
        RECT 27.345 42.715 29.345 42.885 ;
        RECT 30.075 42.195 30.245 52.045 ;
        RECT 30.975 51.355 32.975 51.525 ;
        RECT 33.265 51.355 35.265 51.525 ;
        RECT 35.555 51.355 37.555 51.525 ;
        RECT 37.845 51.355 39.845 51.525 ;
        RECT 40.135 51.355 42.135 51.525 ;
        RECT 42.425 51.355 44.425 51.525 ;
        RECT 44.715 51.355 46.715 51.525 ;
        RECT 47.005 51.355 49.005 51.525 ;
        RECT 30.745 43.100 30.915 51.140 ;
        RECT 33.035 43.100 33.205 51.140 ;
        RECT 35.325 43.100 35.495 51.140 ;
        RECT 37.615 43.100 37.785 51.140 ;
        RECT 39.905 43.100 40.075 51.140 ;
        RECT 42.195 43.100 42.365 51.140 ;
        RECT 44.485 43.100 44.655 51.140 ;
        RECT 46.775 43.100 46.945 51.140 ;
        RECT 49.065 43.100 49.235 51.140 ;
        RECT 30.975 42.715 32.975 42.885 ;
        RECT 33.265 42.715 35.265 42.885 ;
        RECT 35.555 42.715 37.555 42.885 ;
        RECT 37.845 42.715 39.845 42.885 ;
        RECT 40.135 42.715 42.135 42.885 ;
        RECT 42.425 42.715 44.425 42.885 ;
        RECT 44.715 42.715 46.715 42.885 ;
        RECT 47.005 42.715 49.005 42.885 ;
        RECT 49.735 42.195 49.905 52.045 ;
        RECT 50.635 51.355 52.635 51.525 ;
        RECT 52.925 51.355 54.925 51.525 ;
        RECT 55.215 51.355 57.215 51.525 ;
        RECT 57.505 51.355 59.505 51.525 ;
        RECT 59.795 51.355 61.795 51.525 ;
        RECT 62.085 51.355 64.085 51.525 ;
        RECT 64.375 51.355 66.375 51.525 ;
        RECT 66.665 51.355 68.665 51.525 ;
        RECT 50.405 43.100 50.575 51.140 ;
        RECT 52.695 43.100 52.865 51.140 ;
        RECT 54.985 43.100 55.155 51.140 ;
        RECT 57.275 43.100 57.445 51.140 ;
        RECT 59.565 43.100 59.735 51.140 ;
        RECT 61.855 43.100 62.025 51.140 ;
        RECT 64.145 43.100 64.315 51.140 ;
        RECT 66.435 43.100 66.605 51.140 ;
        RECT 68.725 43.100 68.895 51.140 ;
        RECT 50.635 42.715 52.635 42.885 ;
        RECT 52.925 42.715 54.925 42.885 ;
        RECT 55.215 42.715 57.215 42.885 ;
        RECT 57.505 42.715 59.505 42.885 ;
        RECT 59.795 42.715 61.795 42.885 ;
        RECT 62.085 42.715 64.085 42.885 ;
        RECT 64.375 42.715 66.375 42.885 ;
        RECT 66.665 42.715 68.665 42.885 ;
        RECT 69.395 42.195 69.565 52.045 ;
        RECT 70.295 51.355 72.295 51.525 ;
        RECT 72.585 51.355 74.585 51.525 ;
        RECT 74.875 51.355 76.875 51.525 ;
        RECT 77.165 51.355 79.165 51.525 ;
        RECT 79.455 51.355 81.455 51.525 ;
        RECT 81.745 51.355 83.745 51.525 ;
        RECT 84.035 51.355 86.035 51.525 ;
        RECT 86.325 51.355 88.325 51.525 ;
        RECT 70.065 43.100 70.235 51.140 ;
        RECT 72.355 43.100 72.525 51.140 ;
        RECT 74.645 43.100 74.815 51.140 ;
        RECT 76.935 43.100 77.105 51.140 ;
        RECT 79.225 43.100 79.395 51.140 ;
        RECT 81.515 43.100 81.685 51.140 ;
        RECT 83.805 43.100 83.975 51.140 ;
        RECT 86.095 43.100 86.265 51.140 ;
        RECT 88.385 43.100 88.555 51.140 ;
        RECT 70.295 42.715 72.295 42.885 ;
        RECT 72.585 42.715 74.585 42.885 ;
        RECT 74.875 42.715 76.875 42.885 ;
        RECT 77.165 42.715 79.165 42.885 ;
        RECT 79.455 42.715 81.455 42.885 ;
        RECT 81.745 42.715 83.745 42.885 ;
        RECT 84.035 42.715 86.035 42.885 ;
        RECT 86.325 42.715 88.325 42.885 ;
        RECT 89.055 42.195 89.225 52.045 ;
        RECT 89.955 51.355 91.955 51.525 ;
        RECT 92.245 51.355 94.245 51.525 ;
        RECT 94.535 51.355 96.535 51.525 ;
        RECT 96.825 51.355 98.825 51.525 ;
        RECT 99.115 51.355 101.115 51.525 ;
        RECT 101.405 51.355 103.405 51.525 ;
        RECT 103.695 51.355 105.695 51.525 ;
        RECT 105.985 51.355 107.985 51.525 ;
        RECT 89.725 43.100 89.895 51.140 ;
        RECT 92.015 43.100 92.185 51.140 ;
        RECT 94.305 43.100 94.475 51.140 ;
        RECT 96.595 43.100 96.765 51.140 ;
        RECT 98.885 43.100 99.055 51.140 ;
        RECT 101.175 43.100 101.345 51.140 ;
        RECT 103.465 43.100 103.635 51.140 ;
        RECT 105.755 43.100 105.925 51.140 ;
        RECT 108.045 43.100 108.215 51.140 ;
        RECT 89.955 42.715 91.955 42.885 ;
        RECT 92.245 42.715 94.245 42.885 ;
        RECT 94.535 42.715 96.535 42.885 ;
        RECT 96.825 42.715 98.825 42.885 ;
        RECT 99.115 42.715 101.115 42.885 ;
        RECT 101.405 42.715 103.405 42.885 ;
        RECT 103.695 42.715 105.695 42.885 ;
        RECT 105.985 42.715 107.985 42.885 ;
        RECT 108.715 42.195 108.885 52.045 ;
        RECT 109.615 51.355 111.615 51.525 ;
        RECT 111.905 51.355 113.905 51.525 ;
        RECT 114.195 51.355 116.195 51.525 ;
        RECT 116.485 51.355 118.485 51.525 ;
        RECT 118.775 51.355 120.775 51.525 ;
        RECT 121.065 51.355 123.065 51.525 ;
        RECT 123.355 51.355 125.355 51.525 ;
        RECT 125.645 51.355 127.645 51.525 ;
        RECT 109.385 43.100 109.555 51.140 ;
        RECT 111.675 43.100 111.845 51.140 ;
        RECT 113.965 43.100 114.135 51.140 ;
        RECT 116.255 43.100 116.425 51.140 ;
        RECT 118.545 43.100 118.715 51.140 ;
        RECT 120.835 43.100 121.005 51.140 ;
        RECT 123.125 43.100 123.295 51.140 ;
        RECT 125.415 43.100 125.585 51.140 ;
        RECT 127.705 43.100 127.875 51.140 ;
        RECT 109.615 42.715 111.615 42.885 ;
        RECT 111.905 42.715 113.905 42.885 ;
        RECT 114.195 42.715 116.195 42.885 ;
        RECT 116.485 42.715 118.485 42.885 ;
        RECT 118.775 42.715 120.775 42.885 ;
        RECT 121.065 42.715 123.065 42.885 ;
        RECT 123.355 42.715 125.355 42.885 ;
        RECT 125.645 42.715 127.645 42.885 ;
        RECT 128.375 42.195 128.905 52.045 ;
        RECT 10.055 41.665 128.905 42.195 ;
        RECT 10.055 39.070 74.665 39.600 ;
        RECT 10.055 29.310 10.585 39.070 ;
        RECT 11.375 38.380 13.375 38.550 ;
        RECT 13.665 38.380 15.665 38.550 ;
        RECT 15.955 38.380 17.955 38.550 ;
        RECT 18.245 38.380 20.245 38.550 ;
        RECT 11.145 30.170 11.315 38.210 ;
        RECT 13.435 30.170 13.605 38.210 ;
        RECT 15.725 30.170 15.895 38.210 ;
        RECT 18.015 30.170 18.185 38.210 ;
        RECT 20.305 30.170 20.475 38.210 ;
        RECT 11.375 29.830 13.375 30.000 ;
        RECT 13.665 29.830 15.665 30.000 ;
        RECT 15.955 29.830 17.955 30.000 ;
        RECT 18.245 29.830 20.245 30.000 ;
        RECT 21.035 29.310 21.205 39.070 ;
        RECT 21.995 38.380 23.995 38.550 ;
        RECT 24.285 38.380 26.285 38.550 ;
        RECT 26.575 38.380 28.575 38.550 ;
        RECT 28.865 38.380 30.865 38.550 ;
        RECT 21.765 30.170 21.935 38.210 ;
        RECT 24.055 30.170 24.225 38.210 ;
        RECT 26.345 30.170 26.515 38.210 ;
        RECT 28.635 30.170 28.805 38.210 ;
        RECT 30.925 30.170 31.095 38.210 ;
        RECT 21.995 29.830 23.995 30.000 ;
        RECT 24.285 29.830 26.285 30.000 ;
        RECT 26.575 29.830 28.575 30.000 ;
        RECT 28.865 29.830 30.865 30.000 ;
        RECT 31.655 29.310 31.825 39.070 ;
        RECT 32.615 38.380 34.615 38.550 ;
        RECT 34.905 38.380 36.905 38.550 ;
        RECT 37.195 38.380 39.195 38.550 ;
        RECT 39.485 38.380 41.485 38.550 ;
        RECT 32.385 30.170 32.555 38.210 ;
        RECT 34.675 30.170 34.845 38.210 ;
        RECT 36.965 30.170 37.135 38.210 ;
        RECT 39.255 30.170 39.425 38.210 ;
        RECT 41.545 30.170 41.715 38.210 ;
        RECT 32.615 29.830 34.615 30.000 ;
        RECT 34.905 29.830 36.905 30.000 ;
        RECT 37.195 29.830 39.195 30.000 ;
        RECT 39.485 29.830 41.485 30.000 ;
        RECT 42.275 29.310 42.445 39.070 ;
        RECT 43.235 38.380 45.235 38.550 ;
        RECT 45.525 38.380 47.525 38.550 ;
        RECT 47.815 38.380 49.815 38.550 ;
        RECT 50.105 38.380 52.105 38.550 ;
        RECT 43.005 30.170 43.175 38.210 ;
        RECT 45.295 30.170 45.465 38.210 ;
        RECT 47.585 30.170 47.755 38.210 ;
        RECT 49.875 30.170 50.045 38.210 ;
        RECT 52.165 30.170 52.335 38.210 ;
        RECT 43.235 29.830 45.235 30.000 ;
        RECT 45.525 29.830 47.525 30.000 ;
        RECT 47.815 29.830 49.815 30.000 ;
        RECT 50.105 29.830 52.105 30.000 ;
        RECT 52.895 29.310 53.065 39.070 ;
        RECT 53.855 38.380 55.855 38.550 ;
        RECT 56.145 38.380 58.145 38.550 ;
        RECT 58.435 38.380 60.435 38.550 ;
        RECT 60.725 38.380 62.725 38.550 ;
        RECT 53.625 30.170 53.795 38.210 ;
        RECT 55.915 30.170 56.085 38.210 ;
        RECT 58.205 30.170 58.375 38.210 ;
        RECT 60.495 30.170 60.665 38.210 ;
        RECT 62.785 30.170 62.955 38.210 ;
        RECT 53.855 29.830 55.855 30.000 ;
        RECT 56.145 29.830 58.145 30.000 ;
        RECT 58.435 29.830 60.435 30.000 ;
        RECT 60.725 29.830 62.725 30.000 ;
        RECT 63.515 29.310 63.685 39.070 ;
        RECT 64.475 38.380 66.475 38.550 ;
        RECT 66.765 38.380 68.765 38.550 ;
        RECT 69.055 38.380 71.055 38.550 ;
        RECT 71.345 38.380 73.345 38.550 ;
        RECT 64.245 30.170 64.415 38.210 ;
        RECT 66.535 30.170 66.705 38.210 ;
        RECT 68.825 30.170 68.995 38.210 ;
        RECT 71.115 30.170 71.285 38.210 ;
        RECT 73.405 30.170 73.575 38.210 ;
        RECT 64.475 29.830 66.475 30.000 ;
        RECT 66.765 29.830 68.765 30.000 ;
        RECT 69.055 29.830 71.055 30.000 ;
        RECT 71.345 29.830 73.345 30.000 ;
        RECT 74.135 29.310 74.665 39.070 ;
        RECT 10.055 29.140 74.665 29.310 ;
        RECT 10.055 19.380 10.585 29.140 ;
        RECT 11.375 28.450 13.375 28.620 ;
        RECT 13.665 28.450 15.665 28.620 ;
        RECT 15.955 28.450 17.955 28.620 ;
        RECT 18.245 28.450 20.245 28.620 ;
        RECT 11.145 20.240 11.315 28.280 ;
        RECT 13.435 20.240 13.605 28.280 ;
        RECT 15.725 20.240 15.895 28.280 ;
        RECT 18.015 20.240 18.185 28.280 ;
        RECT 20.305 20.240 20.475 28.280 ;
        RECT 11.375 19.900 13.375 20.070 ;
        RECT 13.665 19.900 15.665 20.070 ;
        RECT 15.955 19.900 17.955 20.070 ;
        RECT 18.245 19.900 20.245 20.070 ;
        RECT 21.035 19.380 21.205 29.140 ;
        RECT 21.995 28.450 23.995 28.620 ;
        RECT 24.285 28.450 26.285 28.620 ;
        RECT 26.575 28.450 28.575 28.620 ;
        RECT 28.865 28.450 30.865 28.620 ;
        RECT 21.765 20.240 21.935 28.280 ;
        RECT 24.055 20.240 24.225 28.280 ;
        RECT 26.345 20.240 26.515 28.280 ;
        RECT 28.635 20.240 28.805 28.280 ;
        RECT 30.925 20.240 31.095 28.280 ;
        RECT 21.995 19.900 23.995 20.070 ;
        RECT 24.285 19.900 26.285 20.070 ;
        RECT 26.575 19.900 28.575 20.070 ;
        RECT 28.865 19.900 30.865 20.070 ;
        RECT 31.655 19.380 31.825 29.140 ;
        RECT 32.615 28.450 34.615 28.620 ;
        RECT 34.905 28.450 36.905 28.620 ;
        RECT 37.195 28.450 39.195 28.620 ;
        RECT 39.485 28.450 41.485 28.620 ;
        RECT 32.385 20.240 32.555 28.280 ;
        RECT 34.675 20.240 34.845 28.280 ;
        RECT 36.965 20.240 37.135 28.280 ;
        RECT 39.255 20.240 39.425 28.280 ;
        RECT 41.545 20.240 41.715 28.280 ;
        RECT 32.615 19.900 34.615 20.070 ;
        RECT 34.905 19.900 36.905 20.070 ;
        RECT 37.195 19.900 39.195 20.070 ;
        RECT 39.485 19.900 41.485 20.070 ;
        RECT 42.275 19.380 42.445 29.140 ;
        RECT 43.235 28.450 45.235 28.620 ;
        RECT 45.525 28.450 47.525 28.620 ;
        RECT 47.815 28.450 49.815 28.620 ;
        RECT 50.105 28.450 52.105 28.620 ;
        RECT 43.005 20.240 43.175 28.280 ;
        RECT 45.295 20.240 45.465 28.280 ;
        RECT 47.585 20.240 47.755 28.280 ;
        RECT 49.875 20.240 50.045 28.280 ;
        RECT 52.165 20.240 52.335 28.280 ;
        RECT 43.235 19.900 45.235 20.070 ;
        RECT 45.525 19.900 47.525 20.070 ;
        RECT 47.815 19.900 49.815 20.070 ;
        RECT 50.105 19.900 52.105 20.070 ;
        RECT 52.895 19.380 53.065 29.140 ;
        RECT 53.855 28.450 55.855 28.620 ;
        RECT 56.145 28.450 58.145 28.620 ;
        RECT 58.435 28.450 60.435 28.620 ;
        RECT 60.725 28.450 62.725 28.620 ;
        RECT 53.625 20.240 53.795 28.280 ;
        RECT 55.915 20.240 56.085 28.280 ;
        RECT 58.205 20.240 58.375 28.280 ;
        RECT 60.495 20.240 60.665 28.280 ;
        RECT 62.785 20.240 62.955 28.280 ;
        RECT 53.855 19.900 55.855 20.070 ;
        RECT 56.145 19.900 58.145 20.070 ;
        RECT 58.435 19.900 60.435 20.070 ;
        RECT 60.725 19.900 62.725 20.070 ;
        RECT 63.515 19.380 63.685 29.140 ;
        RECT 64.475 28.450 66.475 28.620 ;
        RECT 66.765 28.450 68.765 28.620 ;
        RECT 69.055 28.450 71.055 28.620 ;
        RECT 71.345 28.450 73.345 28.620 ;
        RECT 64.245 20.240 64.415 28.280 ;
        RECT 66.535 20.240 66.705 28.280 ;
        RECT 68.825 20.240 68.995 28.280 ;
        RECT 71.115 20.240 71.285 28.280 ;
        RECT 73.405 20.240 73.575 28.280 ;
        RECT 64.475 19.900 66.475 20.070 ;
        RECT 66.765 19.900 68.765 20.070 ;
        RECT 69.055 19.900 71.055 20.070 ;
        RECT 71.345 19.900 73.345 20.070 ;
        RECT 74.135 19.380 74.665 29.140 ;
        RECT 10.055 19.210 74.665 19.380 ;
        RECT 10.055 9.450 10.585 19.210 ;
        RECT 11.375 18.520 13.375 18.690 ;
        RECT 13.665 18.520 15.665 18.690 ;
        RECT 15.955 18.520 17.955 18.690 ;
        RECT 18.245 18.520 20.245 18.690 ;
        RECT 11.145 10.310 11.315 18.350 ;
        RECT 13.435 10.310 13.605 18.350 ;
        RECT 15.725 10.310 15.895 18.350 ;
        RECT 18.015 10.310 18.185 18.350 ;
        RECT 20.305 10.310 20.475 18.350 ;
        RECT 11.375 9.970 13.375 10.140 ;
        RECT 13.665 9.970 15.665 10.140 ;
        RECT 15.955 9.970 17.955 10.140 ;
        RECT 18.245 9.970 20.245 10.140 ;
        RECT 21.035 9.450 21.205 19.210 ;
        RECT 21.995 18.520 23.995 18.690 ;
        RECT 24.285 18.520 26.285 18.690 ;
        RECT 26.575 18.520 28.575 18.690 ;
        RECT 28.865 18.520 30.865 18.690 ;
        RECT 21.765 10.310 21.935 18.350 ;
        RECT 24.055 10.310 24.225 18.350 ;
        RECT 26.345 10.310 26.515 18.350 ;
        RECT 28.635 10.310 28.805 18.350 ;
        RECT 30.925 10.310 31.095 18.350 ;
        RECT 21.995 9.970 23.995 10.140 ;
        RECT 24.285 9.970 26.285 10.140 ;
        RECT 26.575 9.970 28.575 10.140 ;
        RECT 28.865 9.970 30.865 10.140 ;
        RECT 31.655 9.450 31.825 19.210 ;
        RECT 32.615 18.520 34.615 18.690 ;
        RECT 34.905 18.520 36.905 18.690 ;
        RECT 37.195 18.520 39.195 18.690 ;
        RECT 39.485 18.520 41.485 18.690 ;
        RECT 32.385 10.310 32.555 18.350 ;
        RECT 34.675 10.310 34.845 18.350 ;
        RECT 36.965 10.310 37.135 18.350 ;
        RECT 39.255 10.310 39.425 18.350 ;
        RECT 41.545 10.310 41.715 18.350 ;
        RECT 32.615 9.970 34.615 10.140 ;
        RECT 34.905 9.970 36.905 10.140 ;
        RECT 37.195 9.970 39.195 10.140 ;
        RECT 39.485 9.970 41.485 10.140 ;
        RECT 42.275 9.450 42.445 19.210 ;
        RECT 43.235 18.520 45.235 18.690 ;
        RECT 45.525 18.520 47.525 18.690 ;
        RECT 47.815 18.520 49.815 18.690 ;
        RECT 50.105 18.520 52.105 18.690 ;
        RECT 43.005 10.310 43.175 18.350 ;
        RECT 45.295 10.310 45.465 18.350 ;
        RECT 47.585 10.310 47.755 18.350 ;
        RECT 49.875 10.310 50.045 18.350 ;
        RECT 52.165 10.310 52.335 18.350 ;
        RECT 43.235 9.970 45.235 10.140 ;
        RECT 45.525 9.970 47.525 10.140 ;
        RECT 47.815 9.970 49.815 10.140 ;
        RECT 50.105 9.970 52.105 10.140 ;
        RECT 52.895 9.450 53.065 19.210 ;
        RECT 53.855 18.520 55.855 18.690 ;
        RECT 56.145 18.520 58.145 18.690 ;
        RECT 58.435 18.520 60.435 18.690 ;
        RECT 60.725 18.520 62.725 18.690 ;
        RECT 53.625 10.310 53.795 18.350 ;
        RECT 55.915 10.310 56.085 18.350 ;
        RECT 58.205 10.310 58.375 18.350 ;
        RECT 60.495 10.310 60.665 18.350 ;
        RECT 62.785 10.310 62.955 18.350 ;
        RECT 53.855 9.970 55.855 10.140 ;
        RECT 56.145 9.970 58.145 10.140 ;
        RECT 58.435 9.970 60.435 10.140 ;
        RECT 60.725 9.970 62.725 10.140 ;
        RECT 63.515 9.450 63.685 19.210 ;
        RECT 64.475 18.520 66.475 18.690 ;
        RECT 66.765 18.520 68.765 18.690 ;
        RECT 69.055 18.520 71.055 18.690 ;
        RECT 71.345 18.520 73.345 18.690 ;
        RECT 64.245 10.310 64.415 18.350 ;
        RECT 66.535 10.310 66.705 18.350 ;
        RECT 68.825 10.310 68.995 18.350 ;
        RECT 71.115 10.310 71.285 18.350 ;
        RECT 73.405 10.310 73.575 18.350 ;
        RECT 64.475 9.970 66.475 10.140 ;
        RECT 66.765 9.970 68.765 10.140 ;
        RECT 69.055 9.970 71.055 10.140 ;
        RECT 71.345 9.970 73.345 10.140 ;
        RECT 74.135 9.450 74.665 19.210 ;
        RECT 10.055 8.920 74.665 9.450 ;
        RECT 79.695 39.070 128.905 39.600 ;
        RECT 79.695 29.310 80.225 39.070 ;
        RECT 80.785 38.210 85.535 39.070 ;
        RECT 80.785 30.170 80.955 38.210 ;
        RECT 83.075 30.170 83.245 38.210 ;
        RECT 85.365 30.170 85.535 38.210 ;
        RECT 81.015 29.830 83.015 30.000 ;
        RECT 83.305 29.830 85.305 30.000 ;
        RECT 86.095 29.310 86.265 39.070 ;
        RECT 87.055 38.380 89.055 38.550 ;
        RECT 89.345 38.380 91.345 38.550 ;
        RECT 86.825 30.170 86.995 38.210 ;
        RECT 89.115 30.170 89.285 38.210 ;
        RECT 91.405 30.170 91.575 38.210 ;
        RECT 87.055 29.830 89.055 30.000 ;
        RECT 89.345 29.830 91.345 30.000 ;
        RECT 92.135 29.310 92.305 39.070 ;
        RECT 93.095 38.380 95.095 38.550 ;
        RECT 95.385 38.380 97.385 38.550 ;
        RECT 92.865 30.170 93.035 38.210 ;
        RECT 95.155 30.170 95.325 38.210 ;
        RECT 97.445 30.170 97.615 38.210 ;
        RECT 93.095 29.830 95.095 30.000 ;
        RECT 95.385 29.830 97.385 30.000 ;
        RECT 98.175 29.310 98.345 39.070 ;
        RECT 99.135 38.380 101.135 38.550 ;
        RECT 101.425 38.380 103.425 38.550 ;
        RECT 98.905 30.170 99.075 38.210 ;
        RECT 101.195 30.170 101.365 38.210 ;
        RECT 103.485 30.170 103.655 38.210 ;
        RECT 99.135 29.830 101.135 30.000 ;
        RECT 101.425 29.830 103.425 30.000 ;
        RECT 104.215 29.310 104.385 39.070 ;
        RECT 105.175 38.380 107.175 38.550 ;
        RECT 107.465 38.380 109.465 38.550 ;
        RECT 104.945 30.170 105.115 38.210 ;
        RECT 107.235 30.170 107.405 38.210 ;
        RECT 109.525 30.170 109.695 38.210 ;
        RECT 105.175 29.830 107.175 30.000 ;
        RECT 107.465 29.830 109.465 30.000 ;
        RECT 110.255 29.310 110.425 39.070 ;
        RECT 111.215 38.380 113.215 38.550 ;
        RECT 113.505 38.380 115.505 38.550 ;
        RECT 110.985 30.170 111.155 38.210 ;
        RECT 113.275 30.170 113.445 38.210 ;
        RECT 115.565 30.170 115.735 38.210 ;
        RECT 111.215 29.830 113.215 30.000 ;
        RECT 113.505 29.830 115.505 30.000 ;
        RECT 116.295 29.310 116.465 39.070 ;
        RECT 117.255 38.380 119.255 38.550 ;
        RECT 119.545 38.380 121.545 38.550 ;
        RECT 117.025 30.170 117.195 38.210 ;
        RECT 119.315 30.170 119.485 38.210 ;
        RECT 121.605 30.170 121.775 38.210 ;
        RECT 117.255 29.830 119.255 30.000 ;
        RECT 119.545 29.830 121.545 30.000 ;
        RECT 122.335 29.310 122.505 39.070 ;
        RECT 123.065 38.210 127.815 39.070 ;
        RECT 123.065 30.170 123.235 38.210 ;
        RECT 125.355 30.170 125.525 38.210 ;
        RECT 127.645 30.170 127.815 38.210 ;
        RECT 123.295 29.830 125.295 30.000 ;
        RECT 125.585 29.830 127.585 30.000 ;
        RECT 128.375 29.310 128.905 39.070 ;
        RECT 79.695 29.140 128.905 29.310 ;
        RECT 79.695 19.380 80.225 29.140 ;
        RECT 81.015 28.450 83.015 28.620 ;
        RECT 83.305 28.450 85.305 28.620 ;
        RECT 80.785 20.240 80.955 28.280 ;
        RECT 83.075 20.240 83.245 28.280 ;
        RECT 85.365 20.240 85.535 28.280 ;
        RECT 80.785 19.380 85.535 20.240 ;
        RECT 86.095 19.380 86.265 29.140 ;
        RECT 87.055 28.450 89.055 28.620 ;
        RECT 89.345 28.450 91.345 28.620 ;
        RECT 86.825 20.240 86.995 28.280 ;
        RECT 89.115 20.240 89.285 28.280 ;
        RECT 91.405 20.240 91.575 28.280 ;
        RECT 87.055 19.900 89.055 20.070 ;
        RECT 89.345 19.900 91.345 20.070 ;
        RECT 92.135 19.380 92.305 29.140 ;
        RECT 93.095 28.450 95.095 28.620 ;
        RECT 95.385 28.450 97.385 28.620 ;
        RECT 92.865 20.240 93.035 28.280 ;
        RECT 95.155 20.240 95.325 28.280 ;
        RECT 97.445 20.240 97.615 28.280 ;
        RECT 93.095 19.900 95.095 20.070 ;
        RECT 95.385 19.900 97.385 20.070 ;
        RECT 98.175 19.380 98.345 29.140 ;
        RECT 99.135 28.450 101.135 28.620 ;
        RECT 101.425 28.450 103.425 28.620 ;
        RECT 98.905 20.240 99.075 28.280 ;
        RECT 101.195 20.240 101.365 28.280 ;
        RECT 103.485 20.240 103.655 28.280 ;
        RECT 99.135 19.900 101.135 20.070 ;
        RECT 101.425 19.900 103.425 20.070 ;
        RECT 104.215 19.380 104.385 29.140 ;
        RECT 105.175 28.450 107.175 28.620 ;
        RECT 107.465 28.450 109.465 28.620 ;
        RECT 104.945 20.240 105.115 28.280 ;
        RECT 107.235 20.240 107.405 28.280 ;
        RECT 109.525 20.240 109.695 28.280 ;
        RECT 105.175 19.900 107.175 20.070 ;
        RECT 107.465 19.900 109.465 20.070 ;
        RECT 110.255 19.380 110.425 29.140 ;
        RECT 111.215 28.450 113.215 28.620 ;
        RECT 113.505 28.450 115.505 28.620 ;
        RECT 110.985 20.240 111.155 28.280 ;
        RECT 113.275 20.240 113.445 28.280 ;
        RECT 115.565 20.240 115.735 28.280 ;
        RECT 111.215 19.900 113.215 20.070 ;
        RECT 113.505 19.900 115.505 20.070 ;
        RECT 116.295 19.380 116.465 29.140 ;
        RECT 117.255 28.450 119.255 28.620 ;
        RECT 119.545 28.450 121.545 28.620 ;
        RECT 117.025 20.240 117.195 28.280 ;
        RECT 119.315 20.240 119.485 28.280 ;
        RECT 121.605 20.240 121.775 28.280 ;
        RECT 117.255 19.900 119.255 20.070 ;
        RECT 119.545 19.900 121.545 20.070 ;
        RECT 122.335 19.380 122.505 29.140 ;
        RECT 123.295 28.450 125.295 28.620 ;
        RECT 125.585 28.450 127.585 28.620 ;
        RECT 123.065 20.240 123.235 28.280 ;
        RECT 125.355 20.240 125.525 28.280 ;
        RECT 127.645 20.240 127.815 28.280 ;
        RECT 123.065 19.380 127.815 20.240 ;
        RECT 128.375 19.380 128.905 29.140 ;
        RECT 79.695 19.210 128.905 19.380 ;
        RECT 79.695 9.450 80.225 19.210 ;
        RECT 81.015 18.520 83.015 18.690 ;
        RECT 83.305 18.520 85.305 18.690 ;
        RECT 80.785 10.310 80.955 18.350 ;
        RECT 83.075 10.310 83.245 18.350 ;
        RECT 85.365 10.310 85.535 18.350 ;
        RECT 80.785 9.450 85.535 10.310 ;
        RECT 86.095 9.450 86.265 19.210 ;
        RECT 87.055 18.520 89.055 18.690 ;
        RECT 89.345 18.520 91.345 18.690 ;
        RECT 86.825 10.310 86.995 18.350 ;
        RECT 89.115 10.310 89.285 18.350 ;
        RECT 91.405 10.310 91.575 18.350 ;
        RECT 86.825 9.450 91.575 10.310 ;
        RECT 92.135 9.450 92.305 19.210 ;
        RECT 93.095 18.520 95.095 18.690 ;
        RECT 95.385 18.520 97.385 18.690 ;
        RECT 92.865 10.310 93.035 18.350 ;
        RECT 95.155 10.310 95.325 18.350 ;
        RECT 97.445 10.310 97.615 18.350 ;
        RECT 92.865 9.450 97.615 10.310 ;
        RECT 98.175 9.450 98.345 19.210 ;
        RECT 99.135 18.520 101.135 18.690 ;
        RECT 101.425 18.520 103.425 18.690 ;
        RECT 98.905 10.310 99.075 18.350 ;
        RECT 101.195 10.310 101.365 18.350 ;
        RECT 103.485 10.310 103.655 18.350 ;
        RECT 98.905 9.450 103.655 10.310 ;
        RECT 104.215 9.450 104.385 19.210 ;
        RECT 105.175 18.520 107.175 18.690 ;
        RECT 107.465 18.520 109.465 18.690 ;
        RECT 104.945 10.310 105.115 18.350 ;
        RECT 107.235 10.310 107.405 18.350 ;
        RECT 109.525 10.310 109.695 18.350 ;
        RECT 104.945 9.450 109.695 10.310 ;
        RECT 110.255 9.450 110.425 19.210 ;
        RECT 111.215 18.520 113.215 18.690 ;
        RECT 113.505 18.520 115.505 18.690 ;
        RECT 110.985 10.310 111.155 18.350 ;
        RECT 113.275 10.310 113.445 18.350 ;
        RECT 115.565 10.310 115.735 18.350 ;
        RECT 110.985 9.450 115.735 10.310 ;
        RECT 116.295 9.450 116.465 19.210 ;
        RECT 117.255 18.520 119.255 18.690 ;
        RECT 119.545 18.520 121.545 18.690 ;
        RECT 117.025 10.310 117.195 18.350 ;
        RECT 119.315 10.310 119.485 18.350 ;
        RECT 121.605 10.310 121.775 18.350 ;
        RECT 117.025 9.450 121.775 10.310 ;
        RECT 122.335 9.450 122.505 19.210 ;
        RECT 123.295 18.520 125.295 18.690 ;
        RECT 125.585 18.520 127.585 18.690 ;
        RECT 123.065 10.310 123.235 18.350 ;
        RECT 125.355 10.310 125.525 18.350 ;
        RECT 127.645 10.310 127.815 18.350 ;
        RECT 123.065 9.450 127.815 10.310 ;
        RECT 128.375 9.450 128.905 19.210 ;
        RECT 135.150 18.895 135.680 104.785 ;
        RECT 136.265 103.615 138.425 104.305 ;
        RECT 136.265 102.445 138.425 103.135 ;
        RECT 136.265 101.275 138.425 101.965 ;
        RECT 136.265 100.105 138.425 100.795 ;
        RECT 136.265 98.935 138.425 99.625 ;
        RECT 136.265 97.765 138.425 98.455 ;
        RECT 136.265 96.595 138.425 97.285 ;
        RECT 136.265 95.425 138.425 96.115 ;
        RECT 136.265 94.255 138.425 94.945 ;
        RECT 136.265 93.085 138.425 93.775 ;
        RECT 136.265 91.915 138.425 92.605 ;
        RECT 136.265 90.745 138.425 91.435 ;
        RECT 136.265 89.575 138.425 90.265 ;
        RECT 136.265 88.405 138.425 89.095 ;
        RECT 136.265 87.235 138.425 87.925 ;
        RECT 136.265 86.065 138.425 86.755 ;
        RECT 136.265 84.895 138.425 85.585 ;
        RECT 136.265 83.725 138.425 84.415 ;
        RECT 136.265 82.555 138.425 83.245 ;
        RECT 136.265 81.385 138.425 82.075 ;
        RECT 136.265 80.215 138.425 80.905 ;
        RECT 136.265 79.045 138.425 79.735 ;
        RECT 136.265 77.875 138.425 78.565 ;
        RECT 136.265 76.705 138.425 77.395 ;
        RECT 136.265 75.535 138.425 76.225 ;
        RECT 136.265 74.365 138.425 75.055 ;
        RECT 136.265 73.195 138.425 73.885 ;
        RECT 136.265 72.025 138.425 72.715 ;
        RECT 136.265 70.855 138.425 71.545 ;
        RECT 136.265 69.685 138.425 70.375 ;
        RECT 136.265 68.515 138.425 69.205 ;
        RECT 136.265 67.345 138.425 68.035 ;
        RECT 136.265 66.175 138.425 66.865 ;
        RECT 136.265 65.005 138.425 65.695 ;
        RECT 136.265 63.835 138.425 64.525 ;
        RECT 136.265 62.665 138.425 63.355 ;
        RECT 136.265 61.495 138.425 62.185 ;
        RECT 136.265 60.325 138.425 61.015 ;
        RECT 136.265 59.155 138.425 59.845 ;
        RECT 136.265 57.985 138.425 58.675 ;
        RECT 136.265 56.815 138.425 57.505 ;
        RECT 136.265 55.645 138.425 56.335 ;
        RECT 136.265 54.475 138.425 55.165 ;
        RECT 136.265 53.305 138.425 53.995 ;
        RECT 136.265 52.135 138.425 52.825 ;
        RECT 136.265 50.965 138.425 51.655 ;
        RECT 136.265 49.795 138.425 50.485 ;
        RECT 136.265 48.625 138.425 49.315 ;
        RECT 136.265 47.455 138.425 48.145 ;
        RECT 136.265 46.285 138.425 46.975 ;
        RECT 136.265 45.115 138.425 45.805 ;
        RECT 136.265 43.945 138.425 44.635 ;
        RECT 136.265 42.775 138.425 43.465 ;
        RECT 136.265 41.605 138.425 42.295 ;
        RECT 136.265 40.435 138.425 41.125 ;
        RECT 136.265 39.265 138.425 39.955 ;
        RECT 136.265 38.095 138.425 38.785 ;
        RECT 136.265 36.925 138.425 37.615 ;
        RECT 136.265 35.755 138.425 36.445 ;
        RECT 136.265 34.585 138.425 35.275 ;
        RECT 136.265 33.415 138.425 34.105 ;
        RECT 136.265 32.245 138.425 32.935 ;
        RECT 136.265 31.075 138.425 31.765 ;
        RECT 136.265 29.905 138.425 30.595 ;
        RECT 136.265 28.735 138.425 29.425 ;
        RECT 136.265 27.565 138.425 28.255 ;
        RECT 136.265 26.395 138.425 27.085 ;
        RECT 136.265 25.225 138.425 25.915 ;
        RECT 136.265 24.055 138.425 24.745 ;
        RECT 136.265 22.885 138.425 23.575 ;
        RECT 136.265 21.715 138.425 22.405 ;
        RECT 136.265 20.545 138.425 21.235 ;
        RECT 136.265 19.375 138.425 20.065 ;
        RECT 139.150 18.895 145.540 104.785 ;
        RECT 146.265 103.615 148.425 104.305 ;
        RECT 146.265 102.445 148.425 103.135 ;
        RECT 146.265 101.275 148.425 101.965 ;
        RECT 146.265 100.105 148.425 100.795 ;
        RECT 146.265 98.935 148.425 99.625 ;
        RECT 146.265 97.765 148.425 98.455 ;
        RECT 146.265 96.595 148.425 97.285 ;
        RECT 146.265 95.425 148.425 96.115 ;
        RECT 146.265 94.255 148.425 94.945 ;
        RECT 146.265 93.085 148.425 93.775 ;
        RECT 146.265 91.915 148.425 92.605 ;
        RECT 146.265 90.745 148.425 91.435 ;
        RECT 146.265 89.575 148.425 90.265 ;
        RECT 146.265 88.405 148.425 89.095 ;
        RECT 146.265 87.235 148.425 87.925 ;
        RECT 146.265 86.065 148.425 86.755 ;
        RECT 146.265 84.895 148.425 85.585 ;
        RECT 146.265 83.725 148.425 84.415 ;
        RECT 146.265 82.555 148.425 83.245 ;
        RECT 146.265 81.385 148.425 82.075 ;
        RECT 146.265 80.215 148.425 80.905 ;
        RECT 146.265 79.045 148.425 79.735 ;
        RECT 146.265 77.875 148.425 78.565 ;
        RECT 146.265 76.705 148.425 77.395 ;
        RECT 146.265 75.535 148.425 76.225 ;
        RECT 146.265 74.365 148.425 75.055 ;
        RECT 146.265 73.195 148.425 73.885 ;
        RECT 146.265 72.025 148.425 72.715 ;
        RECT 146.265 70.855 148.425 71.545 ;
        RECT 146.265 69.685 148.425 70.375 ;
        RECT 146.265 68.515 148.425 69.205 ;
        RECT 146.265 67.345 148.425 68.035 ;
        RECT 146.265 66.175 148.425 66.865 ;
        RECT 146.265 65.005 148.425 65.695 ;
        RECT 146.265 63.835 148.425 64.525 ;
        RECT 146.265 62.665 148.425 63.355 ;
        RECT 146.265 61.495 148.425 62.185 ;
        RECT 146.265 60.325 148.425 61.015 ;
        RECT 146.265 59.155 148.425 59.845 ;
        RECT 146.265 57.985 148.425 58.675 ;
        RECT 146.265 56.815 148.425 57.505 ;
        RECT 146.265 55.645 148.425 56.335 ;
        RECT 146.265 54.475 148.425 55.165 ;
        RECT 146.265 53.305 148.425 53.995 ;
        RECT 146.265 52.135 148.425 52.825 ;
        RECT 146.265 50.965 148.425 51.655 ;
        RECT 146.265 49.795 148.425 50.485 ;
        RECT 146.265 48.625 148.425 49.315 ;
        RECT 146.265 47.455 148.425 48.145 ;
        RECT 146.265 46.285 148.425 46.975 ;
        RECT 146.265 45.115 148.425 45.805 ;
        RECT 146.265 43.945 148.425 44.635 ;
        RECT 146.265 42.775 148.425 43.465 ;
        RECT 146.265 41.605 148.425 42.295 ;
        RECT 146.265 40.435 148.425 41.125 ;
        RECT 146.265 39.265 148.425 39.955 ;
        RECT 146.265 38.095 148.425 38.785 ;
        RECT 146.265 36.925 148.425 37.615 ;
        RECT 146.265 35.755 148.425 36.445 ;
        RECT 146.265 34.585 148.425 35.275 ;
        RECT 146.265 33.415 148.425 34.105 ;
        RECT 146.265 32.245 148.425 32.935 ;
        RECT 146.265 31.075 148.425 31.765 ;
        RECT 146.265 29.905 148.425 30.595 ;
        RECT 146.265 28.735 148.425 29.425 ;
        RECT 146.265 27.565 148.425 28.255 ;
        RECT 146.265 26.395 148.425 27.085 ;
        RECT 146.265 25.225 148.425 25.915 ;
        RECT 146.265 24.055 148.425 24.745 ;
        RECT 146.265 22.885 148.425 23.575 ;
        RECT 146.265 21.715 148.425 22.405 ;
        RECT 146.265 20.545 148.425 21.235 ;
        RECT 146.265 19.375 148.425 20.065 ;
        RECT 149.010 18.895 149.540 104.785 ;
        RECT 135.150 13.490 149.540 18.895 ;
        RECT 79.695 8.920 128.905 9.450 ;
        RECT 155.300 4.700 155.700 180.620 ;
        RECT 165.235 179.815 166.445 180.905 ;
        RECT 166.615 180.955 166.785 181.865 ;
        RECT 167.570 181.795 167.775 182.195 ;
        RECT 167.945 181.965 168.280 182.365 ;
        RECT 168.515 182.000 168.685 182.025 ;
        RECT 166.955 181.125 167.315 181.705 ;
        RECT 167.570 181.625 168.255 181.795 ;
        RECT 167.495 180.955 167.745 181.455 ;
        RECT 166.615 180.785 167.745 180.955 ;
        RECT 166.615 180.015 166.885 180.785 ;
        RECT 167.915 180.595 168.255 181.625 ;
        RECT 167.055 179.815 167.385 180.595 ;
        RECT 167.590 180.420 168.255 180.595 ;
        RECT 168.455 181.625 168.815 182.000 ;
        RECT 169.080 181.625 169.250 182.365 ;
        RECT 169.530 181.795 169.700 182.000 ;
        RECT 169.530 181.625 170.070 181.795 ;
        RECT 168.455 180.970 168.710 181.625 ;
        RECT 168.880 181.125 169.230 181.455 ;
        RECT 169.400 181.125 169.730 181.455 ;
        RECT 167.590 180.015 167.775 180.420 ;
        RECT 167.945 179.815 168.280 180.240 ;
        RECT 168.455 179.985 168.795 180.970 ;
        RECT 168.965 180.585 169.230 181.125 ;
        RECT 169.900 180.925 170.070 181.625 ;
        RECT 169.445 180.755 170.070 180.925 ;
        RECT 170.240 180.995 170.410 182.195 ;
        RECT 170.640 181.715 170.970 182.195 ;
        RECT 171.140 181.895 171.310 182.365 ;
        RECT 171.480 181.715 171.810 182.180 ;
        RECT 170.640 181.545 171.810 181.715 ;
        RECT 172.140 181.625 172.395 182.195 ;
        RECT 172.565 181.965 172.895 182.365 ;
        RECT 173.320 181.830 173.850 182.195 ;
        RECT 174.040 182.025 174.315 182.195 ;
        RECT 174.035 181.855 174.315 182.025 ;
        RECT 173.320 181.795 173.495 181.830 ;
        RECT 172.565 181.625 173.495 181.795 ;
        RECT 170.580 181.165 171.150 181.375 ;
        RECT 171.320 181.165 171.965 181.375 ;
        RECT 170.240 180.585 170.945 180.995 ;
        RECT 172.140 180.955 172.310 181.625 ;
        RECT 172.565 181.455 172.735 181.625 ;
        RECT 172.480 181.125 172.735 181.455 ;
        RECT 172.960 181.125 173.155 181.455 ;
        RECT 168.965 180.415 170.945 180.585 ;
        RECT 168.965 179.815 169.375 180.245 ;
        RECT 170.120 179.815 170.450 180.235 ;
        RECT 170.620 179.985 170.945 180.415 ;
        RECT 171.420 179.815 171.750 180.915 ;
        RECT 172.140 179.985 172.475 180.955 ;
        RECT 172.645 179.815 172.815 180.955 ;
        RECT 172.985 180.155 173.155 181.125 ;
        RECT 173.325 180.495 173.495 181.625 ;
        RECT 173.665 180.835 173.835 181.635 ;
        RECT 174.040 181.035 174.315 181.855 ;
        RECT 174.485 180.835 174.675 182.195 ;
        RECT 174.855 181.830 175.365 182.365 ;
        RECT 175.585 181.555 175.830 182.160 ;
        RECT 176.825 181.815 176.995 182.195 ;
        RECT 177.175 181.985 177.505 182.365 ;
        RECT 176.825 181.645 177.490 181.815 ;
        RECT 177.685 181.690 177.945 182.195 ;
        RECT 174.875 181.385 176.105 181.555 ;
        RECT 173.665 180.665 174.675 180.835 ;
        RECT 174.845 180.820 175.595 181.010 ;
        RECT 173.325 180.325 174.450 180.495 ;
        RECT 174.845 180.155 175.015 180.820 ;
        RECT 175.765 180.575 176.105 181.385 ;
        RECT 176.755 181.095 177.085 181.465 ;
        RECT 177.320 181.390 177.490 181.645 ;
        RECT 177.320 181.060 177.605 181.390 ;
        RECT 177.320 180.915 177.490 181.060 ;
        RECT 172.985 179.985 175.015 180.155 ;
        RECT 175.185 179.815 175.355 180.575 ;
        RECT 175.590 180.165 176.105 180.575 ;
        RECT 176.825 180.745 177.490 180.915 ;
        RECT 177.775 180.890 177.945 181.690 ;
        RECT 178.270 181.715 178.600 182.180 ;
        RECT 178.770 181.895 178.940 182.365 ;
        RECT 179.110 181.715 179.440 182.195 ;
        RECT 178.270 181.545 179.440 181.715 ;
        RECT 178.115 181.165 178.760 181.375 ;
        RECT 178.930 181.165 179.500 181.375 ;
        RECT 179.670 180.995 179.840 182.195 ;
        RECT 180.380 181.795 180.550 182.000 ;
        RECT 176.825 179.985 176.995 180.745 ;
        RECT 177.175 179.815 177.505 180.575 ;
        RECT 177.675 179.985 177.945 180.890 ;
        RECT 178.330 179.815 178.660 180.915 ;
        RECT 179.135 180.585 179.840 180.995 ;
        RECT 180.010 181.625 180.550 181.795 ;
        RECT 180.830 181.625 181.000 182.365 ;
        RECT 181.265 181.625 181.625 182.000 ;
        RECT 180.010 180.925 180.180 181.625 ;
        RECT 180.350 181.125 180.680 181.455 ;
        RECT 180.850 181.125 181.200 181.455 ;
        RECT 180.010 180.755 180.635 180.925 ;
        RECT 180.850 180.585 181.115 181.125 ;
        RECT 181.370 180.970 181.625 181.625 ;
        RECT 181.950 181.715 182.280 182.180 ;
        RECT 182.450 181.895 182.620 182.365 ;
        RECT 182.790 181.715 183.120 182.195 ;
        RECT 181.950 181.545 183.120 181.715 ;
        RECT 181.795 181.165 182.440 181.375 ;
        RECT 182.610 181.165 183.180 181.375 ;
        RECT 183.350 180.995 183.520 182.195 ;
        RECT 184.060 181.795 184.230 182.000 ;
        RECT 179.135 180.415 181.115 180.585 ;
        RECT 179.135 179.985 179.460 180.415 ;
        RECT 179.630 179.815 179.960 180.235 ;
        RECT 180.705 179.815 181.115 180.245 ;
        RECT 181.285 179.985 181.625 180.970 ;
        RECT 182.010 179.815 182.340 180.915 ;
        RECT 182.815 180.585 183.520 180.995 ;
        RECT 183.690 181.625 184.230 181.795 ;
        RECT 184.510 181.625 184.680 182.365 ;
        RECT 184.945 181.625 185.305 182.000 ;
        RECT 185.565 181.815 185.735 182.195 ;
        RECT 185.915 181.985 186.245 182.365 ;
        RECT 185.565 181.645 186.230 181.815 ;
        RECT 186.425 181.690 186.685 182.195 ;
        RECT 183.690 180.925 183.860 181.625 ;
        RECT 184.030 181.125 184.360 181.455 ;
        RECT 184.530 181.125 184.880 181.455 ;
        RECT 183.690 180.755 184.315 180.925 ;
        RECT 184.530 180.585 184.795 181.125 ;
        RECT 185.050 180.970 185.305 181.625 ;
        RECT 185.495 181.095 185.825 181.465 ;
        RECT 186.060 181.390 186.230 181.645 ;
        RECT 182.815 180.415 184.795 180.585 ;
        RECT 182.815 179.985 183.140 180.415 ;
        RECT 183.310 179.815 183.640 180.235 ;
        RECT 184.385 179.815 184.795 180.245 ;
        RECT 184.965 179.985 185.305 180.970 ;
        RECT 186.060 181.060 186.345 181.390 ;
        RECT 186.060 180.915 186.230 181.060 ;
        RECT 185.565 180.745 186.230 180.915 ;
        RECT 186.515 180.890 186.685 181.690 ;
        RECT 185.565 179.985 185.735 180.745 ;
        RECT 185.915 179.815 186.245 180.575 ;
        RECT 186.415 179.985 186.685 180.890 ;
        RECT 186.860 181.625 187.115 182.195 ;
        RECT 187.285 181.965 187.615 182.365 ;
        RECT 188.040 181.830 188.570 182.195 ;
        RECT 188.760 182.025 189.035 182.195 ;
        RECT 188.755 181.855 189.035 182.025 ;
        RECT 188.040 181.795 188.215 181.830 ;
        RECT 187.285 181.625 188.215 181.795 ;
        RECT 186.860 180.955 187.030 181.625 ;
        RECT 187.285 181.455 187.455 181.625 ;
        RECT 187.200 181.125 187.455 181.455 ;
        RECT 187.680 181.125 187.875 181.455 ;
        RECT 186.860 179.985 187.195 180.955 ;
        RECT 187.365 179.815 187.535 180.955 ;
        RECT 187.705 180.155 187.875 181.125 ;
        RECT 188.045 180.495 188.215 181.625 ;
        RECT 188.385 180.835 188.555 181.635 ;
        RECT 188.760 181.035 189.035 181.855 ;
        RECT 189.205 180.835 189.395 182.195 ;
        RECT 189.575 181.830 190.085 182.365 ;
        RECT 190.305 181.555 190.550 182.160 ;
        RECT 190.995 181.640 191.285 182.365 ;
        RECT 192.380 181.715 192.650 181.925 ;
        RECT 192.870 181.905 193.200 182.365 ;
        RECT 193.710 181.905 194.460 182.195 ;
        RECT 189.595 181.385 190.825 181.555 ;
        RECT 192.380 181.545 193.715 181.715 ;
        RECT 188.385 180.665 189.395 180.835 ;
        RECT 189.565 180.820 190.315 181.010 ;
        RECT 188.045 180.325 189.170 180.495 ;
        RECT 189.565 180.155 189.735 180.820 ;
        RECT 190.485 180.575 190.825 181.385 ;
        RECT 193.545 181.375 193.715 181.545 ;
        RECT 192.380 181.135 192.730 181.375 ;
        RECT 192.900 181.135 193.375 181.375 ;
        RECT 193.545 181.125 193.920 181.375 ;
        RECT 187.705 179.985 189.735 180.155 ;
        RECT 189.905 179.815 190.075 180.575 ;
        RECT 190.310 180.165 190.825 180.575 ;
        RECT 190.995 179.815 191.285 180.980 ;
        RECT 193.545 180.955 193.715 181.125 ;
        RECT 192.380 180.785 193.715 180.955 ;
        RECT 192.380 180.625 192.660 180.785 ;
        RECT 194.090 180.615 194.460 181.905 ;
        RECT 192.870 179.815 193.120 180.615 ;
        RECT 193.290 180.445 194.460 180.615 ;
        RECT 194.680 181.625 194.935 182.195 ;
        RECT 195.105 181.965 195.435 182.365 ;
        RECT 195.860 181.830 196.390 182.195 ;
        RECT 195.860 181.795 196.035 181.830 ;
        RECT 195.105 181.625 196.035 181.795 ;
        RECT 194.680 180.955 194.850 181.625 ;
        RECT 195.105 181.455 195.275 181.625 ;
        RECT 195.020 181.125 195.275 181.455 ;
        RECT 195.500 181.125 195.695 181.455 ;
        RECT 193.290 179.985 193.620 180.445 ;
        RECT 193.790 179.815 194.005 180.275 ;
        RECT 194.680 179.985 195.015 180.955 ;
        RECT 195.185 179.815 195.355 180.955 ;
        RECT 195.525 180.155 195.695 181.125 ;
        RECT 195.865 180.495 196.035 181.625 ;
        RECT 196.205 180.835 196.375 181.635 ;
        RECT 196.580 181.345 196.855 182.195 ;
        RECT 196.575 181.175 196.855 181.345 ;
        RECT 196.580 181.035 196.855 181.175 ;
        RECT 197.025 180.835 197.215 182.195 ;
        RECT 197.395 181.830 197.905 182.365 ;
        RECT 198.125 181.555 198.370 182.160 ;
        RECT 198.820 181.625 199.075 182.195 ;
        RECT 199.245 181.965 199.575 182.365 ;
        RECT 200.000 181.830 200.530 182.195 ;
        RECT 200.720 182.025 200.995 182.195 ;
        RECT 200.715 181.855 200.995 182.025 ;
        RECT 200.000 181.795 200.175 181.830 ;
        RECT 199.245 181.625 200.175 181.795 ;
        RECT 197.415 181.385 198.645 181.555 ;
        RECT 196.205 180.665 197.215 180.835 ;
        RECT 197.385 180.820 198.135 181.010 ;
        RECT 195.865 180.325 196.990 180.495 ;
        RECT 197.385 180.155 197.555 180.820 ;
        RECT 198.305 180.575 198.645 181.385 ;
        RECT 195.525 179.985 197.555 180.155 ;
        RECT 197.725 179.815 197.895 180.575 ;
        RECT 198.130 180.165 198.645 180.575 ;
        RECT 198.820 180.955 198.990 181.625 ;
        RECT 199.245 181.455 199.415 181.625 ;
        RECT 199.160 181.125 199.415 181.455 ;
        RECT 199.640 181.125 199.835 181.455 ;
        RECT 198.820 179.985 199.155 180.955 ;
        RECT 199.325 179.815 199.495 180.955 ;
        RECT 199.665 180.155 199.835 181.125 ;
        RECT 200.005 180.495 200.175 181.625 ;
        RECT 200.345 180.835 200.515 181.635 ;
        RECT 200.720 181.035 200.995 181.855 ;
        RECT 201.165 180.835 201.355 182.195 ;
        RECT 201.535 181.830 202.045 182.365 ;
        RECT 202.265 181.555 202.510 182.160 ;
        RECT 203.045 181.815 203.215 182.195 ;
        RECT 203.395 181.985 203.725 182.365 ;
        RECT 203.045 181.645 203.710 181.815 ;
        RECT 203.905 181.690 204.165 182.195 ;
        RECT 201.555 181.385 202.785 181.555 ;
        RECT 200.345 180.665 201.355 180.835 ;
        RECT 201.525 180.820 202.275 181.010 ;
        RECT 200.005 180.325 201.130 180.495 ;
        RECT 201.525 180.155 201.695 180.820 ;
        RECT 202.445 180.575 202.785 181.385 ;
        RECT 202.975 181.095 203.305 181.465 ;
        RECT 203.540 181.390 203.710 181.645 ;
        RECT 203.540 181.060 203.825 181.390 ;
        RECT 203.540 180.915 203.710 181.060 ;
        RECT 199.665 179.985 201.695 180.155 ;
        RECT 201.865 179.815 202.035 180.575 ;
        RECT 202.270 180.165 202.785 180.575 ;
        RECT 203.045 180.745 203.710 180.915 ;
        RECT 203.995 180.890 204.165 181.690 ;
        RECT 204.425 181.815 204.595 182.195 ;
        RECT 204.775 181.985 205.105 182.365 ;
        RECT 204.425 181.645 205.090 181.815 ;
        RECT 205.285 181.690 205.545 182.195 ;
        RECT 204.355 181.095 204.685 181.465 ;
        RECT 204.920 181.390 205.090 181.645 ;
        RECT 204.920 181.060 205.205 181.390 ;
        RECT 204.920 180.915 205.090 181.060 ;
        RECT 203.045 179.985 203.215 180.745 ;
        RECT 203.395 179.815 203.725 180.575 ;
        RECT 203.895 179.985 204.165 180.890 ;
        RECT 204.425 180.745 205.090 180.915 ;
        RECT 205.375 180.890 205.545 181.690 ;
        RECT 205.805 181.815 205.975 182.195 ;
        RECT 206.155 181.985 206.485 182.365 ;
        RECT 205.805 181.645 206.470 181.815 ;
        RECT 206.665 181.690 206.925 182.195 ;
        RECT 205.735 181.095 206.065 181.465 ;
        RECT 206.300 181.390 206.470 181.645 ;
        RECT 206.300 181.060 206.585 181.390 ;
        RECT 206.300 180.915 206.470 181.060 ;
        RECT 204.425 179.985 204.595 180.745 ;
        RECT 204.775 179.815 205.105 180.575 ;
        RECT 205.275 179.985 205.545 180.890 ;
        RECT 205.805 180.745 206.470 180.915 ;
        RECT 206.755 180.890 206.925 181.690 ;
        RECT 207.185 181.815 207.355 182.190 ;
        RECT 207.525 181.985 207.855 182.365 ;
        RECT 208.025 182.025 209.100 182.195 ;
        RECT 208.025 181.815 208.195 182.025 ;
        RECT 207.185 181.645 208.195 181.815 ;
        RECT 208.420 181.685 208.760 181.855 ;
        RECT 208.930 181.690 209.100 182.025 ;
        RECT 208.420 181.515 208.710 181.685 ;
        RECT 207.160 181.005 207.505 181.455 ;
        RECT 205.805 179.985 205.975 180.745 ;
        RECT 206.155 179.815 206.485 180.575 ;
        RECT 206.655 179.985 206.925 180.890 ;
        RECT 207.155 180.835 207.505 181.005 ;
        RECT 207.815 180.835 208.250 181.455 ;
        RECT 208.420 180.995 208.590 181.515 ;
        RECT 209.270 181.345 209.630 182.020 ;
        RECT 209.810 181.645 210.100 182.365 ;
        RECT 210.390 182.025 211.990 182.195 ;
        RECT 210.390 181.655 210.560 182.025 ;
        RECT 211.635 181.985 211.990 182.025 ;
        RECT 212.160 181.905 212.330 182.365 ;
        RECT 210.730 181.605 211.060 181.855 ;
        RECT 210.745 181.530 211.060 181.605 ;
        RECT 211.230 181.735 211.400 181.855 ;
        RECT 212.505 181.735 212.750 182.155 ;
        RECT 213.020 181.985 213.350 182.365 ;
        RECT 213.520 181.795 213.695 182.125 ;
        RECT 214.040 182.035 214.210 182.195 ;
        RECT 214.040 181.865 214.570 182.035 ;
        RECT 214.740 182.025 215.735 182.195 ;
        RECT 214.740 181.865 214.910 182.025 ;
        RECT 211.230 181.565 212.750 181.735 ;
        RECT 209.090 181.165 209.630 181.345 ;
        RECT 209.270 181.055 209.630 181.165 ;
        RECT 208.420 180.825 209.055 180.995 ;
        RECT 209.270 180.825 210.075 181.055 ;
        RECT 207.185 180.485 208.715 180.655 ;
        RECT 207.185 179.985 207.355 180.485 ;
        RECT 208.545 180.325 208.715 180.485 ;
        RECT 208.885 180.495 209.055 180.825 ;
        RECT 208.885 180.325 209.215 180.495 ;
        RECT 207.525 179.815 207.855 180.195 ;
        RECT 208.025 180.155 208.195 180.315 ;
        RECT 209.385 180.155 209.555 180.655 ;
        RECT 208.025 179.985 209.555 180.155 ;
        RECT 209.725 179.985 210.075 180.825 ;
        RECT 210.275 180.455 210.575 181.455 ;
        RECT 210.745 181.005 210.915 181.530 ;
        RECT 211.230 181.525 211.400 181.565 ;
        RECT 211.085 181.345 211.415 181.355 ;
        RECT 211.085 181.185 211.470 181.345 ;
        RECT 211.300 181.175 211.470 181.185 ;
        RECT 211.810 181.005 212.055 181.395 ;
        RECT 210.745 180.835 211.505 181.005 ;
        RECT 211.755 180.835 212.055 181.005 ;
        RECT 210.245 179.815 210.575 180.195 ;
        RECT 210.835 180.155 211.005 180.665 ;
        RECT 211.175 180.325 211.505 180.835 ;
        RECT 211.810 180.775 212.055 180.835 ;
        RECT 212.260 180.775 212.590 181.395 ;
        RECT 213.065 180.775 213.355 181.455 ;
        RECT 213.525 181.345 213.695 181.795 ;
        RECT 213.990 181.515 214.230 181.685 ;
        RECT 213.525 181.175 213.815 181.345 ;
        RECT 211.675 180.365 212.740 180.535 ;
        RECT 211.675 180.155 211.845 180.365 ;
        RECT 210.835 179.985 211.845 180.155 ;
        RECT 212.070 179.815 212.400 180.195 ;
        RECT 212.570 179.985 212.740 180.365 ;
        RECT 213.525 180.315 213.695 181.175 ;
        RECT 212.990 179.815 213.340 180.195 ;
        RECT 213.510 179.985 213.695 180.315 ;
        RECT 213.990 180.315 214.160 181.515 ;
        RECT 214.400 180.695 214.570 181.865 ;
        RECT 215.220 181.685 215.395 181.855 ;
        RECT 214.980 181.525 215.395 181.685 ;
        RECT 215.565 181.735 215.735 182.025 ;
        RECT 215.905 181.905 216.075 182.365 ;
        RECT 215.565 181.565 216.135 181.735 ;
        RECT 214.980 181.515 215.390 181.525 ;
        RECT 215.200 181.175 215.655 181.345 ;
        RECT 215.965 180.785 216.135 181.565 ;
        RECT 214.400 180.465 215.185 180.695 ;
        RECT 214.855 180.325 215.185 180.465 ;
        RECT 215.485 180.615 216.135 180.785 ;
        RECT 213.990 179.985 214.200 180.315 ;
        RECT 214.370 180.155 214.700 180.195 ;
        RECT 215.485 180.155 215.655 180.615 ;
        RECT 214.370 179.985 215.655 180.155 ;
        RECT 215.825 179.815 216.155 180.195 ;
        RECT 216.325 179.985 216.585 182.195 ;
        RECT 216.755 181.640 217.045 182.365 ;
        RECT 217.305 181.815 217.475 182.190 ;
        RECT 217.645 181.985 217.975 182.365 ;
        RECT 218.145 182.025 219.220 182.195 ;
        RECT 218.145 181.815 218.315 182.025 ;
        RECT 217.305 181.645 218.315 181.815 ;
        RECT 218.540 181.685 218.880 181.855 ;
        RECT 219.050 181.690 219.220 182.025 ;
        RECT 218.540 181.515 218.830 181.685 ;
        RECT 217.280 181.345 217.625 181.455 ;
        RECT 217.275 181.175 217.625 181.345 ;
        RECT 216.755 179.815 217.045 180.980 ;
        RECT 217.280 180.835 217.625 181.175 ;
        RECT 217.935 180.835 218.370 181.455 ;
        RECT 218.540 180.995 218.710 181.515 ;
        RECT 219.390 181.345 219.750 182.020 ;
        RECT 219.930 181.645 220.220 182.365 ;
        RECT 220.510 182.025 222.110 182.195 ;
        RECT 220.510 181.655 220.680 182.025 ;
        RECT 221.755 181.985 222.110 182.025 ;
        RECT 222.280 181.905 222.450 182.365 ;
        RECT 220.850 181.605 221.180 181.855 ;
        RECT 220.865 181.530 221.180 181.605 ;
        RECT 221.350 181.735 221.520 181.855 ;
        RECT 222.625 181.735 222.870 182.155 ;
        RECT 223.140 181.985 223.470 182.365 ;
        RECT 223.640 181.795 223.815 182.125 ;
        RECT 224.160 182.035 224.330 182.195 ;
        RECT 224.160 181.865 224.690 182.035 ;
        RECT 224.860 182.025 225.855 182.195 ;
        RECT 224.860 181.865 225.030 182.025 ;
        RECT 221.350 181.565 222.870 181.735 ;
        RECT 219.210 181.165 219.750 181.345 ;
        RECT 219.390 181.055 219.750 181.165 ;
        RECT 218.540 180.825 219.175 180.995 ;
        RECT 219.390 180.825 220.195 181.055 ;
        RECT 217.305 180.485 218.835 180.655 ;
        RECT 217.305 179.985 217.475 180.485 ;
        RECT 218.665 180.325 218.835 180.485 ;
        RECT 219.005 180.495 219.175 180.825 ;
        RECT 219.005 180.325 219.335 180.495 ;
        RECT 217.645 179.815 217.975 180.195 ;
        RECT 218.145 180.155 218.315 180.315 ;
        RECT 219.505 180.155 219.675 180.655 ;
        RECT 218.145 179.985 219.675 180.155 ;
        RECT 219.845 179.985 220.195 180.825 ;
        RECT 220.395 180.455 220.695 181.455 ;
        RECT 220.865 181.005 221.035 181.530 ;
        RECT 221.350 181.525 221.520 181.565 ;
        RECT 221.205 181.345 221.535 181.355 ;
        RECT 221.205 181.185 221.590 181.345 ;
        RECT 221.420 181.175 221.590 181.185 ;
        RECT 221.930 181.005 222.175 181.395 ;
        RECT 220.865 180.835 221.625 181.005 ;
        RECT 221.875 180.835 222.175 181.005 ;
        RECT 220.365 179.815 220.695 180.195 ;
        RECT 220.955 180.155 221.125 180.665 ;
        RECT 221.295 180.325 221.625 180.835 ;
        RECT 221.930 180.775 222.175 180.835 ;
        RECT 222.380 180.775 222.710 181.395 ;
        RECT 223.185 180.775 223.475 181.455 ;
        RECT 223.645 181.345 223.815 181.795 ;
        RECT 224.110 181.515 224.350 181.685 ;
        RECT 223.645 181.175 223.935 181.345 ;
        RECT 221.795 180.365 222.860 180.535 ;
        RECT 221.795 180.155 221.965 180.365 ;
        RECT 220.955 179.985 221.965 180.155 ;
        RECT 222.190 179.815 222.520 180.195 ;
        RECT 222.690 179.985 222.860 180.365 ;
        RECT 223.645 180.315 223.815 181.175 ;
        RECT 223.110 179.815 223.460 180.195 ;
        RECT 223.630 179.985 223.815 180.315 ;
        RECT 224.110 180.315 224.280 181.515 ;
        RECT 224.520 180.695 224.690 181.865 ;
        RECT 225.340 181.685 225.515 181.855 ;
        RECT 225.100 181.525 225.515 181.685 ;
        RECT 225.685 181.735 225.855 182.025 ;
        RECT 226.025 181.905 226.195 182.365 ;
        RECT 225.685 181.565 226.255 181.735 ;
        RECT 225.100 181.515 225.510 181.525 ;
        RECT 225.320 181.175 225.775 181.345 ;
        RECT 226.085 180.785 226.255 181.565 ;
        RECT 224.520 180.465 225.305 180.695 ;
        RECT 224.975 180.325 225.305 180.465 ;
        RECT 225.605 180.615 226.255 180.785 ;
        RECT 224.110 179.985 224.320 180.315 ;
        RECT 224.490 180.155 224.820 180.195 ;
        RECT 225.605 180.155 225.775 180.615 ;
        RECT 224.490 179.985 225.775 180.155 ;
        RECT 225.945 179.815 226.275 180.195 ;
        RECT 226.445 179.985 226.705 182.195 ;
        RECT 226.965 181.815 227.135 182.190 ;
        RECT 227.305 181.985 227.635 182.365 ;
        RECT 227.805 182.025 228.880 182.195 ;
        RECT 227.805 181.815 227.975 182.025 ;
        RECT 226.965 181.645 227.975 181.815 ;
        RECT 228.200 181.685 228.540 181.855 ;
        RECT 228.710 181.690 228.880 182.025 ;
        RECT 228.200 181.515 228.490 181.685 ;
        RECT 226.940 181.005 227.285 181.455 ;
        RECT 226.935 180.835 227.285 181.005 ;
        RECT 227.595 180.835 228.030 181.455 ;
        RECT 228.200 180.995 228.370 181.515 ;
        RECT 229.050 181.345 229.410 182.020 ;
        RECT 229.590 181.645 229.880 182.365 ;
        RECT 230.170 182.025 231.770 182.195 ;
        RECT 230.170 181.655 230.340 182.025 ;
        RECT 231.415 181.985 231.770 182.025 ;
        RECT 231.940 181.905 232.110 182.365 ;
        RECT 230.510 181.605 230.840 181.855 ;
        RECT 230.525 181.530 230.840 181.605 ;
        RECT 231.010 181.735 231.180 181.855 ;
        RECT 232.285 181.735 232.530 182.155 ;
        RECT 232.800 181.985 233.130 182.365 ;
        RECT 233.300 181.795 233.475 182.125 ;
        RECT 233.820 182.035 233.990 182.195 ;
        RECT 233.820 181.865 234.350 182.035 ;
        RECT 234.520 182.025 235.515 182.195 ;
        RECT 234.520 181.865 234.690 182.025 ;
        RECT 231.010 181.565 232.530 181.735 ;
        RECT 228.870 181.165 229.410 181.345 ;
        RECT 229.050 181.055 229.410 181.165 ;
        RECT 228.200 180.825 228.835 180.995 ;
        RECT 229.050 180.825 229.855 181.055 ;
        RECT 226.965 180.485 228.495 180.655 ;
        RECT 226.965 179.985 227.135 180.485 ;
        RECT 228.325 180.325 228.495 180.485 ;
        RECT 228.665 180.495 228.835 180.825 ;
        RECT 228.665 180.325 228.995 180.495 ;
        RECT 227.305 179.815 227.635 180.195 ;
        RECT 227.805 180.155 227.975 180.315 ;
        RECT 229.165 180.155 229.335 180.655 ;
        RECT 227.805 179.985 229.335 180.155 ;
        RECT 229.505 179.985 229.855 180.825 ;
        RECT 230.055 180.455 230.355 181.455 ;
        RECT 230.525 181.005 230.695 181.530 ;
        RECT 231.010 181.525 231.180 181.565 ;
        RECT 230.865 181.345 231.195 181.355 ;
        RECT 230.865 181.185 231.250 181.345 ;
        RECT 231.080 181.175 231.250 181.185 ;
        RECT 230.525 180.835 231.285 181.005 ;
        RECT 230.025 179.815 230.355 180.195 ;
        RECT 230.615 180.155 230.785 180.665 ;
        RECT 230.955 180.325 231.285 180.835 ;
        RECT 231.590 180.775 231.835 181.395 ;
        RECT 232.040 181.005 232.370 181.395 ;
        RECT 232.040 180.835 232.395 181.005 ;
        RECT 232.040 180.775 232.370 180.835 ;
        RECT 232.845 180.775 233.135 181.455 ;
        RECT 233.305 181.345 233.475 181.795 ;
        RECT 233.770 181.515 234.010 181.685 ;
        RECT 233.305 181.175 233.595 181.345 ;
        RECT 231.455 180.365 232.520 180.535 ;
        RECT 231.455 180.155 231.625 180.365 ;
        RECT 230.615 179.985 231.625 180.155 ;
        RECT 231.850 179.815 232.180 180.195 ;
        RECT 232.350 179.985 232.520 180.365 ;
        RECT 233.305 180.315 233.475 181.175 ;
        RECT 232.770 179.815 233.120 180.195 ;
        RECT 233.290 179.985 233.475 180.315 ;
        RECT 233.770 180.315 233.940 181.515 ;
        RECT 234.180 180.695 234.350 181.865 ;
        RECT 235.000 181.685 235.175 181.855 ;
        RECT 234.760 181.525 235.175 181.685 ;
        RECT 235.345 181.735 235.515 182.025 ;
        RECT 235.685 181.905 235.855 182.365 ;
        RECT 235.345 181.565 235.915 181.735 ;
        RECT 234.760 181.515 235.170 181.525 ;
        RECT 234.980 181.175 235.435 181.345 ;
        RECT 235.745 180.785 235.915 181.565 ;
        RECT 234.180 180.465 234.965 180.695 ;
        RECT 234.635 180.325 234.965 180.465 ;
        RECT 235.265 180.615 235.915 180.785 ;
        RECT 233.770 179.985 233.980 180.315 ;
        RECT 234.150 180.155 234.480 180.195 ;
        RECT 235.265 180.155 235.435 180.615 ;
        RECT 234.150 179.985 235.435 180.155 ;
        RECT 235.605 179.815 235.935 180.195 ;
        RECT 236.105 179.985 236.365 182.195 ;
        RECT 236.535 181.690 236.795 182.195 ;
        RECT 236.975 181.985 237.305 182.365 ;
        RECT 237.485 181.815 237.655 182.195 ;
        RECT 236.535 180.890 236.705 181.690 ;
        RECT 236.990 181.645 237.655 181.815 ;
        RECT 236.990 181.390 237.160 181.645 ;
        RECT 237.915 181.615 239.125 182.365 ;
        RECT 236.875 181.060 237.160 181.390 ;
        RECT 237.395 181.095 237.725 181.465 ;
        RECT 236.990 180.915 237.160 181.060 ;
        RECT 236.535 179.985 236.805 180.890 ;
        RECT 236.990 180.745 237.655 180.915 ;
        RECT 236.975 179.815 237.305 180.575 ;
        RECT 237.485 179.985 237.655 180.745 ;
        RECT 237.915 180.905 238.435 181.445 ;
        RECT 238.605 181.075 239.125 181.615 ;
        RECT 237.915 179.815 239.125 180.905 ;
        RECT 165.150 179.645 239.210 179.815 ;
        RECT 165.235 178.555 166.445 179.645 ;
        RECT 165.235 177.845 165.755 178.385 ;
        RECT 165.925 178.015 166.445 178.555 ;
        RECT 167.165 178.715 167.335 179.475 ;
        RECT 167.515 178.885 167.845 179.645 ;
        RECT 167.165 178.545 167.830 178.715 ;
        RECT 168.015 178.570 168.285 179.475 ;
        RECT 167.660 178.400 167.830 178.545 ;
        RECT 167.095 177.995 167.425 178.365 ;
        RECT 167.660 178.070 167.945 178.400 ;
        RECT 165.235 177.095 166.445 177.845 ;
        RECT 167.660 177.815 167.830 178.070 ;
        RECT 167.165 177.645 167.830 177.815 ;
        RECT 168.115 177.770 168.285 178.570 ;
        RECT 168.545 178.715 168.715 179.475 ;
        RECT 168.895 178.885 169.225 179.645 ;
        RECT 168.545 178.545 169.210 178.715 ;
        RECT 169.395 178.570 169.665 179.475 ;
        RECT 170.330 178.845 170.580 179.645 ;
        RECT 170.750 179.015 171.080 179.475 ;
        RECT 171.250 179.185 171.465 179.645 ;
        RECT 170.750 178.845 171.920 179.015 ;
        RECT 169.040 178.400 169.210 178.545 ;
        RECT 168.475 177.995 168.805 178.365 ;
        RECT 169.040 178.070 169.325 178.400 ;
        RECT 169.040 177.815 169.210 178.070 ;
        RECT 167.165 177.265 167.335 177.645 ;
        RECT 167.515 177.095 167.845 177.475 ;
        RECT 168.025 177.265 168.285 177.770 ;
        RECT 168.545 177.645 169.210 177.815 ;
        RECT 169.495 177.770 169.665 178.570 ;
        RECT 169.840 178.675 170.120 178.835 ;
        RECT 169.840 178.505 171.175 178.675 ;
        RECT 171.005 178.335 171.175 178.505 ;
        RECT 169.840 178.085 170.190 178.325 ;
        RECT 170.360 178.085 170.835 178.325 ;
        RECT 171.005 178.085 171.380 178.335 ;
        RECT 171.005 177.915 171.175 178.085 ;
        RECT 168.545 177.265 168.715 177.645 ;
        RECT 168.895 177.095 169.225 177.475 ;
        RECT 169.405 177.265 169.665 177.770 ;
        RECT 169.840 177.745 171.175 177.915 ;
        RECT 169.840 177.535 170.110 177.745 ;
        RECT 171.550 177.555 171.920 178.845 ;
        RECT 172.350 178.545 172.680 179.645 ;
        RECT 173.155 179.045 173.480 179.475 ;
        RECT 173.650 179.225 173.980 179.645 ;
        RECT 174.725 179.215 175.135 179.645 ;
        RECT 173.155 178.875 175.135 179.045 ;
        RECT 173.155 178.465 173.860 178.875 ;
        RECT 172.135 178.085 172.780 178.295 ;
        RECT 172.950 178.085 173.520 178.295 ;
        RECT 170.330 177.095 170.660 177.555 ;
        RECT 171.170 177.265 171.920 177.555 ;
        RECT 172.290 177.745 173.460 177.915 ;
        RECT 172.290 177.280 172.620 177.745 ;
        RECT 172.790 177.095 172.960 177.565 ;
        RECT 173.130 177.265 173.460 177.745 ;
        RECT 173.690 177.265 173.860 178.465 ;
        RECT 174.030 178.535 174.655 178.705 ;
        RECT 174.030 177.835 174.200 178.535 ;
        RECT 174.870 178.335 175.135 178.875 ;
        RECT 175.305 178.490 175.645 179.475 ;
        RECT 176.310 178.845 176.560 179.645 ;
        RECT 176.730 179.015 177.060 179.475 ;
        RECT 177.230 179.185 177.445 179.645 ;
        RECT 176.730 178.845 177.900 179.015 ;
        RECT 175.820 178.675 176.100 178.835 ;
        RECT 175.820 178.505 177.155 178.675 ;
        RECT 174.370 178.005 174.700 178.335 ;
        RECT 174.870 178.005 175.220 178.335 ;
        RECT 175.390 177.835 175.645 178.490 ;
        RECT 176.985 178.335 177.155 178.505 ;
        RECT 175.820 178.085 176.170 178.325 ;
        RECT 176.340 178.085 176.815 178.325 ;
        RECT 176.985 178.085 177.360 178.335 ;
        RECT 176.985 177.915 177.155 178.085 ;
        RECT 174.030 177.665 174.570 177.835 ;
        RECT 174.400 177.460 174.570 177.665 ;
        RECT 174.850 177.095 175.020 177.835 ;
        RECT 175.285 177.460 175.645 177.835 ;
        RECT 175.820 177.745 177.155 177.915 ;
        RECT 175.820 177.535 176.090 177.745 ;
        RECT 177.530 177.555 177.900 178.845 ;
        RECT 178.115 178.480 178.405 179.645 ;
        RECT 178.665 178.715 178.835 179.475 ;
        RECT 179.015 178.885 179.345 179.645 ;
        RECT 178.665 178.545 179.330 178.715 ;
        RECT 179.515 178.570 179.785 179.475 ;
        RECT 179.160 178.400 179.330 178.545 ;
        RECT 178.595 177.995 178.925 178.365 ;
        RECT 179.160 178.070 179.445 178.400 ;
        RECT 176.310 177.095 176.640 177.555 ;
        RECT 177.150 177.265 177.900 177.555 ;
        RECT 178.115 177.095 178.405 177.820 ;
        RECT 179.160 177.815 179.330 178.070 ;
        RECT 178.665 177.645 179.330 177.815 ;
        RECT 179.615 177.770 179.785 178.570 ;
        RECT 180.045 178.715 180.215 179.475 ;
        RECT 180.395 178.885 180.725 179.645 ;
        RECT 180.045 178.545 180.710 178.715 ;
        RECT 180.895 178.570 181.165 179.475 ;
        RECT 180.540 178.400 180.710 178.545 ;
        RECT 179.975 177.995 180.305 178.365 ;
        RECT 180.540 178.070 180.825 178.400 ;
        RECT 180.540 177.815 180.710 178.070 ;
        RECT 178.665 177.265 178.835 177.645 ;
        RECT 179.015 177.095 179.345 177.475 ;
        RECT 179.525 177.265 179.785 177.770 ;
        RECT 180.045 177.645 180.710 177.815 ;
        RECT 180.995 177.770 181.165 178.570 ;
        RECT 181.425 178.715 181.595 179.475 ;
        RECT 181.775 178.885 182.105 179.645 ;
        RECT 181.425 178.545 182.090 178.715 ;
        RECT 182.275 178.570 182.545 179.475 ;
        RECT 181.920 178.400 182.090 178.545 ;
        RECT 181.355 177.995 181.685 178.365 ;
        RECT 181.920 178.070 182.205 178.400 ;
        RECT 181.920 177.815 182.090 178.070 ;
        RECT 180.045 177.265 180.215 177.645 ;
        RECT 180.395 177.095 180.725 177.475 ;
        RECT 180.905 177.265 181.165 177.770 ;
        RECT 181.425 177.645 182.090 177.815 ;
        RECT 182.375 177.770 182.545 178.570 ;
        RECT 181.425 177.265 181.595 177.645 ;
        RECT 181.775 177.095 182.105 177.475 ;
        RECT 182.285 177.265 182.545 177.770 ;
        RECT 182.715 178.570 182.985 179.475 ;
        RECT 183.155 178.885 183.485 179.645 ;
        RECT 183.665 178.715 183.835 179.475 ;
        RECT 182.715 177.770 182.885 178.570 ;
        RECT 183.170 178.545 183.835 178.715 ;
        RECT 184.185 178.715 184.355 179.475 ;
        RECT 184.535 178.885 184.865 179.645 ;
        RECT 184.185 178.545 184.850 178.715 ;
        RECT 185.035 178.570 185.305 179.475 ;
        RECT 183.170 178.400 183.340 178.545 ;
        RECT 183.055 178.070 183.340 178.400 ;
        RECT 184.680 178.400 184.850 178.545 ;
        RECT 183.170 177.815 183.340 178.070 ;
        RECT 183.575 177.995 183.905 178.365 ;
        RECT 184.115 177.995 184.445 178.365 ;
        RECT 184.680 178.070 184.965 178.400 ;
        RECT 184.680 177.815 184.850 178.070 ;
        RECT 182.715 177.265 182.975 177.770 ;
        RECT 183.170 177.645 183.835 177.815 ;
        RECT 183.155 177.095 183.485 177.475 ;
        RECT 183.665 177.265 183.835 177.645 ;
        RECT 184.185 177.645 184.850 177.815 ;
        RECT 185.135 177.770 185.305 178.570 ;
        RECT 184.185 177.265 184.355 177.645 ;
        RECT 184.535 177.095 184.865 177.475 ;
        RECT 185.045 177.265 185.305 177.770 ;
        RECT 185.480 178.505 185.815 179.475 ;
        RECT 185.985 178.505 186.155 179.645 ;
        RECT 186.325 179.305 188.355 179.475 ;
        RECT 185.480 177.835 185.650 178.505 ;
        RECT 186.325 178.335 186.495 179.305 ;
        RECT 185.820 178.005 186.075 178.335 ;
        RECT 186.300 178.005 186.495 178.335 ;
        RECT 186.665 178.965 187.790 179.135 ;
        RECT 185.905 177.835 186.075 178.005 ;
        RECT 186.665 177.835 186.835 178.965 ;
        RECT 185.480 177.265 185.735 177.835 ;
        RECT 185.905 177.665 186.835 177.835 ;
        RECT 187.005 178.625 188.015 178.795 ;
        RECT 187.005 177.825 187.175 178.625 ;
        RECT 187.380 178.285 187.655 178.425 ;
        RECT 187.375 178.115 187.655 178.285 ;
        RECT 186.660 177.630 186.835 177.665 ;
        RECT 185.905 177.095 186.235 177.495 ;
        RECT 186.660 177.265 187.190 177.630 ;
        RECT 187.380 177.265 187.655 178.115 ;
        RECT 187.825 177.265 188.015 178.625 ;
        RECT 188.185 178.640 188.355 179.305 ;
        RECT 188.525 178.885 188.695 179.645 ;
        RECT 188.930 178.885 189.445 179.295 ;
        RECT 188.185 178.450 188.935 178.640 ;
        RECT 189.105 178.075 189.445 178.885 ;
        RECT 189.705 178.715 189.875 179.475 ;
        RECT 190.055 178.885 190.385 179.645 ;
        RECT 189.705 178.545 190.370 178.715 ;
        RECT 190.555 178.570 190.825 179.475 ;
        RECT 190.200 178.400 190.370 178.545 ;
        RECT 188.215 177.905 189.445 178.075 ;
        RECT 189.635 177.995 189.965 178.365 ;
        RECT 190.200 178.070 190.485 178.400 ;
        RECT 188.195 177.095 188.705 177.630 ;
        RECT 188.925 177.300 189.170 177.905 ;
        RECT 190.200 177.815 190.370 178.070 ;
        RECT 189.705 177.645 190.370 177.815 ;
        RECT 190.655 177.770 190.825 178.570 ;
        RECT 190.995 178.480 191.285 179.645 ;
        RECT 191.545 178.715 191.715 179.475 ;
        RECT 191.895 178.885 192.225 179.645 ;
        RECT 191.545 178.545 192.210 178.715 ;
        RECT 192.395 178.570 192.665 179.475 ;
        RECT 192.040 178.400 192.210 178.545 ;
        RECT 191.475 177.995 191.805 178.365 ;
        RECT 192.040 178.070 192.325 178.400 ;
        RECT 189.705 177.265 189.875 177.645 ;
        RECT 190.055 177.095 190.385 177.475 ;
        RECT 190.565 177.265 190.825 177.770 ;
        RECT 190.995 177.095 191.285 177.820 ;
        RECT 192.040 177.815 192.210 178.070 ;
        RECT 191.545 177.645 192.210 177.815 ;
        RECT 192.495 177.770 192.665 178.570 ;
        RECT 191.545 177.265 191.715 177.645 ;
        RECT 191.895 177.095 192.225 177.475 ;
        RECT 192.405 177.265 192.665 177.770 ;
        RECT 192.840 178.505 193.175 179.475 ;
        RECT 193.345 178.505 193.515 179.645 ;
        RECT 193.685 179.305 195.715 179.475 ;
        RECT 192.840 177.835 193.010 178.505 ;
        RECT 193.685 178.335 193.855 179.305 ;
        RECT 193.180 178.005 193.435 178.335 ;
        RECT 193.660 178.005 193.855 178.335 ;
        RECT 194.025 178.965 195.150 179.135 ;
        RECT 193.265 177.835 193.435 178.005 ;
        RECT 194.025 177.835 194.195 178.965 ;
        RECT 192.840 177.265 193.095 177.835 ;
        RECT 193.265 177.665 194.195 177.835 ;
        RECT 194.365 178.625 195.375 178.795 ;
        RECT 194.365 177.825 194.535 178.625 ;
        RECT 194.740 178.285 195.015 178.425 ;
        RECT 194.735 178.115 195.015 178.285 ;
        RECT 194.020 177.630 194.195 177.665 ;
        RECT 193.265 177.095 193.595 177.495 ;
        RECT 194.020 177.265 194.550 177.630 ;
        RECT 194.740 177.265 195.015 178.115 ;
        RECT 195.185 177.265 195.375 178.625 ;
        RECT 195.545 178.640 195.715 179.305 ;
        RECT 195.885 178.885 196.055 179.645 ;
        RECT 196.290 178.885 196.805 179.295 ;
        RECT 195.545 178.450 196.295 178.640 ;
        RECT 196.465 178.075 196.805 178.885 ;
        RECT 197.065 178.715 197.235 179.475 ;
        RECT 197.415 178.885 197.745 179.645 ;
        RECT 197.065 178.545 197.730 178.715 ;
        RECT 197.915 178.570 198.185 179.475 ;
        RECT 197.560 178.400 197.730 178.545 ;
        RECT 195.575 177.905 196.805 178.075 ;
        RECT 196.995 177.995 197.325 178.365 ;
        RECT 197.560 178.070 197.845 178.400 ;
        RECT 195.555 177.095 196.065 177.630 ;
        RECT 196.285 177.300 196.530 177.905 ;
        RECT 197.560 177.815 197.730 178.070 ;
        RECT 197.065 177.645 197.730 177.815 ;
        RECT 198.015 177.770 198.185 178.570 ;
        RECT 197.065 177.265 197.235 177.645 ;
        RECT 197.415 177.095 197.745 177.475 ;
        RECT 197.925 177.265 198.185 177.770 ;
        RECT 198.360 178.505 198.695 179.475 ;
        RECT 198.865 178.505 199.035 179.645 ;
        RECT 199.205 179.305 201.235 179.475 ;
        RECT 198.360 177.835 198.530 178.505 ;
        RECT 199.205 178.335 199.375 179.305 ;
        RECT 198.700 178.005 198.955 178.335 ;
        RECT 199.180 178.005 199.375 178.335 ;
        RECT 199.545 178.965 200.670 179.135 ;
        RECT 198.785 177.835 198.955 178.005 ;
        RECT 199.545 177.835 199.715 178.965 ;
        RECT 198.360 177.265 198.615 177.835 ;
        RECT 198.785 177.665 199.715 177.835 ;
        RECT 199.885 178.625 200.895 178.795 ;
        RECT 199.885 177.825 200.055 178.625 ;
        RECT 199.540 177.630 199.715 177.665 ;
        RECT 198.785 177.095 199.115 177.495 ;
        RECT 199.540 177.265 200.070 177.630 ;
        RECT 200.260 177.605 200.535 178.425 ;
        RECT 200.255 177.435 200.535 177.605 ;
        RECT 200.260 177.265 200.535 177.435 ;
        RECT 200.705 177.265 200.895 178.625 ;
        RECT 201.065 178.640 201.235 179.305 ;
        RECT 201.405 178.885 201.575 179.645 ;
        RECT 201.810 178.885 202.325 179.295 ;
        RECT 201.065 178.450 201.815 178.640 ;
        RECT 201.985 178.075 202.325 178.885 ;
        RECT 202.585 178.715 202.755 179.475 ;
        RECT 202.935 178.885 203.265 179.645 ;
        RECT 202.585 178.545 203.250 178.715 ;
        RECT 203.435 178.570 203.705 179.475 ;
        RECT 203.080 178.400 203.250 178.545 ;
        RECT 201.095 177.905 202.325 178.075 ;
        RECT 202.515 177.995 202.845 178.365 ;
        RECT 203.080 178.070 203.365 178.400 ;
        RECT 201.075 177.095 201.585 177.630 ;
        RECT 201.805 177.300 202.050 177.905 ;
        RECT 203.080 177.815 203.250 178.070 ;
        RECT 202.585 177.645 203.250 177.815 ;
        RECT 203.535 177.770 203.705 178.570 ;
        RECT 203.875 178.480 204.165 179.645 ;
        RECT 204.885 178.715 205.055 179.475 ;
        RECT 205.235 178.885 205.565 179.645 ;
        RECT 204.885 178.545 205.550 178.715 ;
        RECT 205.735 178.570 206.005 179.475 ;
        RECT 205.380 178.400 205.550 178.545 ;
        RECT 204.815 177.995 205.145 178.365 ;
        RECT 205.380 178.070 205.665 178.400 ;
        RECT 202.585 177.265 202.755 177.645 ;
        RECT 202.935 177.095 203.265 177.475 ;
        RECT 203.445 177.265 203.705 177.770 ;
        RECT 203.875 177.095 204.165 177.820 ;
        RECT 205.380 177.815 205.550 178.070 ;
        RECT 204.885 177.645 205.550 177.815 ;
        RECT 205.835 177.770 206.005 178.570 ;
        RECT 204.885 177.265 205.055 177.645 ;
        RECT 205.235 177.095 205.565 177.475 ;
        RECT 205.745 177.265 206.005 177.770 ;
        RECT 207.095 177.265 207.355 179.475 ;
        RECT 207.525 179.265 207.855 179.645 ;
        RECT 208.025 179.305 209.310 179.475 ;
        RECT 208.025 178.845 208.195 179.305 ;
        RECT 208.980 179.265 209.310 179.305 ;
        RECT 209.480 179.145 209.690 179.475 ;
        RECT 207.545 178.675 208.195 178.845 ;
        RECT 208.495 178.995 208.825 179.135 ;
        RECT 208.495 178.765 209.280 178.995 ;
        RECT 207.545 177.895 207.715 178.675 ;
        RECT 208.025 178.115 208.480 178.285 ;
        RECT 208.290 177.935 208.700 177.945 ;
        RECT 207.545 177.725 208.115 177.895 ;
        RECT 207.605 177.095 207.775 177.555 ;
        RECT 207.945 177.435 208.115 177.725 ;
        RECT 208.285 177.775 208.700 177.935 ;
        RECT 208.285 177.605 208.460 177.775 ;
        RECT 209.110 177.595 209.280 178.765 ;
        RECT 209.520 177.945 209.690 179.145 ;
        RECT 209.985 179.145 210.170 179.475 ;
        RECT 210.340 179.265 210.690 179.645 ;
        RECT 209.985 178.285 210.155 179.145 ;
        RECT 210.940 179.095 211.110 179.475 ;
        RECT 211.280 179.265 211.610 179.645 ;
        RECT 211.835 179.305 212.845 179.475 ;
        RECT 211.835 179.095 212.005 179.305 ;
        RECT 210.940 178.925 212.005 179.095 ;
        RECT 209.865 178.115 210.155 178.285 ;
        RECT 209.450 177.775 209.690 177.945 ;
        RECT 209.985 177.665 210.155 178.115 ;
        RECT 210.325 178.005 210.615 178.685 ;
        RECT 211.090 178.065 211.420 178.685 ;
        RECT 211.625 178.285 211.870 178.685 ;
        RECT 212.175 178.625 212.505 179.135 ;
        RECT 212.675 178.795 212.845 179.305 ;
        RECT 213.105 179.265 213.435 179.645 ;
        RECT 212.175 178.455 212.935 178.625 ;
        RECT 211.625 178.115 211.925 178.285 ;
        RECT 212.210 178.275 212.380 178.285 ;
        RECT 212.210 178.115 212.595 178.275 ;
        RECT 211.625 178.065 211.870 178.115 ;
        RECT 212.265 178.105 212.595 178.115 ;
        RECT 212.280 177.895 212.450 177.935 ;
        RECT 212.765 177.930 212.935 178.455 ;
        RECT 213.105 178.005 213.405 179.005 ;
        RECT 213.605 178.635 213.955 179.475 ;
        RECT 214.125 179.305 215.655 179.475 ;
        RECT 214.125 178.805 214.295 179.305 ;
        RECT 215.485 179.145 215.655 179.305 ;
        RECT 215.825 179.265 216.155 179.645 ;
        RECT 214.465 178.965 214.795 179.135 ;
        RECT 214.625 178.635 214.795 178.965 ;
        RECT 214.965 178.975 215.135 179.135 ;
        RECT 216.325 178.975 216.495 179.475 ;
        RECT 214.965 178.805 216.495 178.975 ;
        RECT 213.605 178.405 214.410 178.635 ;
        RECT 214.625 178.465 215.260 178.635 ;
        RECT 214.050 178.295 214.410 178.405 ;
        RECT 214.050 178.115 214.590 178.295 ;
        RECT 210.930 177.725 212.450 177.895 ;
        RECT 208.770 177.435 208.940 177.595 ;
        RECT 207.945 177.265 208.940 177.435 ;
        RECT 209.110 177.425 209.640 177.595 ;
        RECT 209.470 177.265 209.640 177.425 ;
        RECT 209.985 177.335 210.160 177.665 ;
        RECT 210.330 177.095 210.660 177.475 ;
        RECT 210.930 177.305 211.175 177.725 ;
        RECT 212.280 177.605 212.450 177.725 ;
        RECT 212.620 177.855 212.935 177.930 ;
        RECT 212.620 177.605 212.950 177.855 ;
        RECT 211.350 177.095 211.520 177.555 ;
        RECT 211.690 177.435 212.045 177.475 ;
        RECT 213.120 177.435 213.290 177.805 ;
        RECT 211.690 177.265 213.290 177.435 ;
        RECT 213.580 177.095 213.870 177.815 ;
        RECT 214.050 177.440 214.410 178.115 ;
        RECT 215.090 177.945 215.260 178.465 ;
        RECT 215.430 178.005 215.865 178.625 ;
        RECT 216.175 178.455 216.525 178.625 ;
        RECT 216.755 178.480 217.045 179.645 ;
        RECT 217.305 178.715 217.475 179.475 ;
        RECT 217.655 178.885 217.985 179.645 ;
        RECT 217.305 178.545 217.970 178.715 ;
        RECT 218.155 178.570 218.425 179.475 ;
        RECT 216.175 178.005 216.520 178.455 ;
        RECT 217.800 178.400 217.970 178.545 ;
        RECT 217.235 177.995 217.565 178.365 ;
        RECT 217.800 178.070 218.085 178.400 ;
        RECT 214.970 177.775 215.260 177.945 ;
        RECT 214.580 177.435 214.750 177.770 ;
        RECT 214.920 177.605 215.260 177.775 ;
        RECT 215.485 177.645 216.495 177.815 ;
        RECT 215.485 177.435 215.655 177.645 ;
        RECT 214.580 177.265 215.655 177.435 ;
        RECT 215.825 177.095 216.155 177.475 ;
        RECT 216.325 177.270 216.495 177.645 ;
        RECT 216.755 177.095 217.045 177.820 ;
        RECT 217.800 177.815 217.970 178.070 ;
        RECT 217.305 177.645 217.970 177.815 ;
        RECT 218.255 177.770 218.425 178.570 ;
        RECT 218.685 178.715 218.855 179.475 ;
        RECT 219.035 178.885 219.365 179.645 ;
        RECT 218.685 178.545 219.350 178.715 ;
        RECT 219.535 178.570 219.805 179.475 ;
        RECT 220.065 178.975 220.235 179.475 ;
        RECT 220.405 179.265 220.735 179.645 ;
        RECT 220.905 179.305 222.435 179.475 ;
        RECT 220.905 179.145 221.075 179.305 ;
        RECT 221.425 178.975 221.595 179.135 ;
        RECT 220.065 178.805 221.595 178.975 ;
        RECT 221.765 178.965 222.095 179.135 ;
        RECT 221.765 178.635 221.935 178.965 ;
        RECT 222.265 178.805 222.435 179.305 ;
        RECT 222.605 178.635 222.955 179.475 ;
        RECT 223.125 179.265 223.455 179.645 ;
        RECT 223.715 179.305 224.725 179.475 ;
        RECT 219.180 178.400 219.350 178.545 ;
        RECT 218.615 177.995 218.945 178.365 ;
        RECT 219.180 178.070 219.465 178.400 ;
        RECT 219.180 177.815 219.350 178.070 ;
        RECT 217.305 177.265 217.475 177.645 ;
        RECT 217.655 177.095 217.985 177.475 ;
        RECT 218.165 177.265 218.425 177.770 ;
        RECT 218.685 177.645 219.350 177.815 ;
        RECT 219.635 177.770 219.805 178.570 ;
        RECT 220.040 178.285 220.385 178.625 ;
        RECT 220.035 178.115 220.385 178.285 ;
        RECT 220.040 178.005 220.385 178.115 ;
        RECT 220.695 178.005 221.130 178.625 ;
        RECT 221.300 178.465 221.935 178.635 ;
        RECT 221.300 177.945 221.470 178.465 ;
        RECT 222.150 178.405 222.955 178.635 ;
        RECT 222.150 178.295 222.510 178.405 ;
        RECT 221.970 178.115 222.510 178.295 ;
        RECT 218.685 177.265 218.855 177.645 ;
        RECT 219.035 177.095 219.365 177.475 ;
        RECT 219.545 177.265 219.805 177.770 ;
        RECT 220.065 177.645 221.075 177.815 ;
        RECT 220.065 177.270 220.235 177.645 ;
        RECT 220.405 177.095 220.735 177.475 ;
        RECT 220.905 177.435 221.075 177.645 ;
        RECT 221.300 177.775 221.590 177.945 ;
        RECT 221.300 177.605 221.640 177.775 ;
        RECT 221.810 177.435 221.980 177.770 ;
        RECT 222.150 177.440 222.510 178.115 ;
        RECT 223.155 178.005 223.455 179.005 ;
        RECT 223.715 178.795 223.885 179.305 ;
        RECT 224.055 178.625 224.385 179.135 ;
        RECT 224.555 179.095 224.725 179.305 ;
        RECT 224.950 179.265 225.280 179.645 ;
        RECT 225.450 179.095 225.620 179.475 ;
        RECT 225.870 179.265 226.220 179.645 ;
        RECT 226.390 179.145 226.575 179.475 ;
        RECT 224.555 178.925 225.620 179.095 ;
        RECT 223.625 178.455 224.385 178.625 ;
        RECT 223.625 177.930 223.795 178.455 ;
        RECT 224.690 178.285 224.935 178.685 ;
        RECT 224.180 178.275 224.350 178.285 ;
        RECT 223.965 178.115 224.350 178.275 ;
        RECT 224.635 178.115 224.935 178.285 ;
        RECT 223.965 178.105 224.295 178.115 ;
        RECT 224.690 178.065 224.935 178.115 ;
        RECT 225.140 178.625 225.470 178.685 ;
        RECT 225.140 178.455 225.495 178.625 ;
        RECT 225.140 178.065 225.470 178.455 ;
        RECT 225.945 178.005 226.235 178.685 ;
        RECT 226.405 178.285 226.575 179.145 ;
        RECT 226.870 179.145 227.080 179.475 ;
        RECT 227.250 179.305 228.535 179.475 ;
        RECT 227.250 179.265 227.580 179.305 ;
        RECT 226.405 178.115 226.695 178.285 ;
        RECT 223.625 177.855 223.940 177.930 ;
        RECT 220.905 177.265 221.980 177.435 ;
        RECT 222.690 177.095 222.980 177.815 ;
        RECT 223.270 177.435 223.440 177.805 ;
        RECT 223.610 177.605 223.940 177.855 ;
        RECT 224.110 177.895 224.280 177.935 ;
        RECT 224.110 177.725 225.630 177.895 ;
        RECT 224.110 177.605 224.280 177.725 ;
        RECT 224.515 177.435 224.870 177.475 ;
        RECT 223.270 177.265 224.870 177.435 ;
        RECT 225.040 177.095 225.210 177.555 ;
        RECT 225.385 177.305 225.630 177.725 ;
        RECT 226.405 177.665 226.575 178.115 ;
        RECT 226.870 177.945 227.040 179.145 ;
        RECT 227.735 178.995 228.065 179.135 ;
        RECT 227.280 178.765 228.065 178.995 ;
        RECT 228.365 178.845 228.535 179.305 ;
        RECT 228.705 179.265 229.035 179.645 ;
        RECT 226.870 177.775 227.110 177.945 ;
        RECT 225.900 177.095 226.230 177.475 ;
        RECT 226.400 177.335 226.575 177.665 ;
        RECT 227.280 177.595 227.450 178.765 ;
        RECT 228.365 178.675 229.015 178.845 ;
        RECT 228.080 178.115 228.535 178.285 ;
        RECT 227.860 177.935 228.270 177.945 ;
        RECT 227.860 177.775 228.275 177.935 ;
        RECT 228.845 177.895 229.015 178.675 ;
        RECT 228.100 177.605 228.275 177.775 ;
        RECT 228.445 177.725 229.015 177.895 ;
        RECT 226.920 177.425 227.450 177.595 ;
        RECT 227.620 177.435 227.790 177.595 ;
        RECT 228.445 177.435 228.615 177.725 ;
        RECT 226.920 177.265 227.090 177.425 ;
        RECT 227.620 177.265 228.615 177.435 ;
        RECT 228.785 177.095 228.955 177.555 ;
        RECT 229.205 177.265 229.465 179.475 ;
        RECT 229.635 178.480 229.925 179.645 ;
        RECT 230.095 178.570 230.365 179.475 ;
        RECT 230.535 178.885 230.865 179.645 ;
        RECT 231.045 178.715 231.215 179.475 ;
        RECT 229.635 177.095 229.925 177.820 ;
        RECT 230.095 177.770 230.265 178.570 ;
        RECT 230.550 178.545 231.215 178.715 ;
        RECT 231.475 178.570 231.745 179.475 ;
        RECT 231.915 178.885 232.245 179.645 ;
        RECT 232.425 178.715 232.595 179.475 ;
        RECT 230.550 178.400 230.720 178.545 ;
        RECT 230.435 178.070 230.720 178.400 ;
        RECT 230.550 177.815 230.720 178.070 ;
        RECT 230.955 177.995 231.285 178.365 ;
        RECT 230.095 177.265 230.355 177.770 ;
        RECT 230.550 177.645 231.215 177.815 ;
        RECT 230.535 177.095 230.865 177.475 ;
        RECT 231.045 177.265 231.215 177.645 ;
        RECT 231.475 177.770 231.645 178.570 ;
        RECT 231.930 178.545 232.595 178.715 ;
        RECT 232.855 178.570 233.125 179.475 ;
        RECT 233.295 178.885 233.625 179.645 ;
        RECT 233.805 178.715 233.975 179.475 ;
        RECT 231.930 178.400 232.100 178.545 ;
        RECT 231.815 178.070 232.100 178.400 ;
        RECT 231.930 177.815 232.100 178.070 ;
        RECT 232.335 177.995 232.665 178.365 ;
        RECT 231.475 177.265 231.735 177.770 ;
        RECT 231.930 177.645 232.595 177.815 ;
        RECT 231.915 177.095 232.245 177.475 ;
        RECT 232.425 177.265 232.595 177.645 ;
        RECT 232.855 177.770 233.025 178.570 ;
        RECT 233.310 178.545 233.975 178.715 ;
        RECT 234.235 178.570 234.505 179.475 ;
        RECT 234.675 178.885 235.005 179.645 ;
        RECT 235.185 178.715 235.355 179.475 ;
        RECT 233.310 178.400 233.480 178.545 ;
        RECT 233.195 178.070 233.480 178.400 ;
        RECT 233.310 177.815 233.480 178.070 ;
        RECT 233.715 177.995 234.045 178.365 ;
        RECT 232.855 177.265 233.115 177.770 ;
        RECT 233.310 177.645 233.975 177.815 ;
        RECT 233.295 177.095 233.625 177.475 ;
        RECT 233.805 177.265 233.975 177.645 ;
        RECT 234.235 177.770 234.405 178.570 ;
        RECT 234.690 178.545 235.355 178.715 ;
        RECT 235.615 178.570 235.885 179.475 ;
        RECT 236.055 178.885 236.385 179.645 ;
        RECT 236.565 178.715 236.735 179.475 ;
        RECT 234.690 178.400 234.860 178.545 ;
        RECT 234.575 178.070 234.860 178.400 ;
        RECT 234.690 177.815 234.860 178.070 ;
        RECT 235.095 177.995 235.425 178.365 ;
        RECT 234.235 177.265 234.495 177.770 ;
        RECT 234.690 177.645 235.355 177.815 ;
        RECT 234.675 177.095 235.005 177.475 ;
        RECT 235.185 177.265 235.355 177.645 ;
        RECT 235.615 177.770 235.785 178.570 ;
        RECT 236.070 178.545 236.735 178.715 ;
        RECT 237.915 178.555 239.125 179.645 ;
        RECT 236.070 178.400 236.240 178.545 ;
        RECT 235.955 178.070 236.240 178.400 ;
        RECT 236.070 177.815 236.240 178.070 ;
        RECT 236.475 177.995 236.805 178.365 ;
        RECT 237.915 178.015 238.435 178.555 ;
        RECT 238.605 177.845 239.125 178.385 ;
        RECT 235.615 177.265 235.875 177.770 ;
        RECT 236.070 177.645 236.735 177.815 ;
        RECT 236.055 177.095 236.385 177.475 ;
        RECT 236.565 177.265 236.735 177.645 ;
        RECT 237.915 177.095 239.125 177.845 ;
        RECT 165.150 176.925 239.210 177.095 ;
        RECT 162.095 106.340 311.135 106.510 ;
        RECT 162.180 105.590 163.390 106.340 ;
        RECT 162.180 105.050 162.700 105.590 ;
        RECT 164.025 105.500 164.285 106.340 ;
        RECT 164.460 105.595 164.715 106.170 ;
        RECT 164.885 105.960 165.215 106.340 ;
        RECT 165.430 105.790 165.600 106.170 ;
        RECT 164.885 105.620 165.600 105.790 ;
        RECT 162.870 104.880 163.390 105.420 ;
        RECT 162.180 103.790 163.390 104.880 ;
        RECT 164.025 103.790 164.285 104.940 ;
        RECT 164.460 104.865 164.630 105.595 ;
        RECT 164.885 105.430 165.055 105.620 ;
        RECT 165.865 105.500 166.125 106.340 ;
        RECT 166.300 105.595 166.555 106.170 ;
        RECT 166.725 105.960 167.055 106.340 ;
        RECT 167.270 105.790 167.440 106.170 ;
        RECT 166.725 105.620 167.440 105.790 ;
        RECT 164.800 105.100 165.055 105.430 ;
        RECT 164.885 104.890 165.055 105.100 ;
        RECT 165.335 105.070 165.690 105.440 ;
        RECT 164.460 103.960 164.715 104.865 ;
        RECT 164.885 104.720 165.600 104.890 ;
        RECT 164.885 103.790 165.215 104.550 ;
        RECT 165.430 103.960 165.600 104.720 ;
        RECT 165.865 103.790 166.125 104.940 ;
        RECT 166.300 104.865 166.470 105.595 ;
        RECT 166.725 105.430 166.895 105.620 ;
        RECT 167.705 105.500 167.965 106.340 ;
        RECT 168.140 105.595 168.395 106.170 ;
        RECT 168.565 105.960 168.895 106.340 ;
        RECT 169.110 105.790 169.280 106.170 ;
        RECT 168.565 105.620 169.280 105.790 ;
        RECT 166.640 105.100 166.895 105.430 ;
        RECT 166.725 104.890 166.895 105.100 ;
        RECT 167.175 105.070 167.530 105.440 ;
        RECT 166.300 103.960 166.555 104.865 ;
        RECT 166.725 104.720 167.440 104.890 ;
        RECT 166.725 103.790 167.055 104.550 ;
        RECT 167.270 103.960 167.440 104.720 ;
        RECT 167.705 103.790 167.965 104.940 ;
        RECT 168.140 104.865 168.310 105.595 ;
        RECT 168.565 105.430 168.735 105.620 ;
        RECT 169.545 105.500 169.805 106.340 ;
        RECT 169.980 105.595 170.235 106.170 ;
        RECT 170.405 105.960 170.735 106.340 ;
        RECT 170.950 105.790 171.120 106.170 ;
        RECT 170.405 105.620 171.120 105.790 ;
        RECT 168.480 105.100 168.735 105.430 ;
        RECT 168.565 104.890 168.735 105.100 ;
        RECT 169.015 105.070 169.370 105.440 ;
        RECT 168.140 103.960 168.395 104.865 ;
        RECT 168.565 104.720 169.280 104.890 ;
        RECT 168.565 103.790 168.895 104.550 ;
        RECT 169.110 103.960 169.280 104.720 ;
        RECT 169.545 103.790 169.805 104.940 ;
        RECT 169.980 104.865 170.150 105.595 ;
        RECT 170.405 105.430 170.575 105.620 ;
        RECT 171.385 105.500 171.645 106.340 ;
        RECT 171.820 105.595 172.075 106.170 ;
        RECT 172.245 105.960 172.575 106.340 ;
        RECT 172.790 105.790 172.960 106.170 ;
        RECT 172.245 105.620 172.960 105.790 ;
        RECT 173.310 105.790 173.480 106.170 ;
        RECT 173.695 105.960 174.025 106.340 ;
        RECT 173.310 105.620 174.025 105.790 ;
        RECT 170.320 105.100 170.575 105.430 ;
        RECT 170.405 104.890 170.575 105.100 ;
        RECT 170.855 105.070 171.210 105.440 ;
        RECT 169.980 103.960 170.235 104.865 ;
        RECT 170.405 104.720 171.120 104.890 ;
        RECT 170.405 103.790 170.735 104.550 ;
        RECT 170.950 103.960 171.120 104.720 ;
        RECT 171.385 103.790 171.645 104.940 ;
        RECT 171.820 104.865 171.990 105.595 ;
        RECT 172.245 105.430 172.415 105.620 ;
        RECT 172.160 105.100 172.415 105.430 ;
        RECT 172.245 104.890 172.415 105.100 ;
        RECT 172.695 105.070 173.050 105.440 ;
        RECT 173.220 105.070 173.575 105.440 ;
        RECT 173.855 105.430 174.025 105.620 ;
        RECT 174.195 105.595 174.450 106.170 ;
        RECT 173.855 105.100 174.110 105.430 ;
        RECT 173.855 104.890 174.025 105.100 ;
        RECT 171.820 103.960 172.075 104.865 ;
        RECT 172.245 104.720 172.960 104.890 ;
        RECT 172.245 103.790 172.575 104.550 ;
        RECT 172.790 103.960 172.960 104.720 ;
        RECT 173.310 104.720 174.025 104.890 ;
        RECT 174.280 104.865 174.450 105.595 ;
        RECT 174.625 105.500 174.885 106.340 ;
        RECT 175.060 105.615 175.350 106.340 ;
        RECT 175.525 105.600 175.780 106.170 ;
        RECT 175.950 105.940 176.280 106.340 ;
        RECT 176.705 105.805 177.235 106.170 ;
        RECT 176.705 105.770 176.880 105.805 ;
        RECT 175.950 105.600 176.880 105.770 ;
        RECT 173.310 103.960 173.480 104.720 ;
        RECT 173.695 103.790 174.025 104.550 ;
        RECT 174.195 103.960 174.450 104.865 ;
        RECT 174.625 103.790 174.885 104.940 ;
        RECT 175.060 103.790 175.350 104.955 ;
        RECT 175.525 104.930 175.695 105.600 ;
        RECT 175.950 105.430 176.120 105.600 ;
        RECT 175.865 105.100 176.120 105.430 ;
        RECT 176.345 105.100 176.540 105.430 ;
        RECT 175.525 103.960 175.860 104.930 ;
        RECT 176.030 103.790 176.200 104.930 ;
        RECT 176.370 104.130 176.540 105.100 ;
        RECT 176.710 104.470 176.880 105.600 ;
        RECT 177.050 104.810 177.220 105.610 ;
        RECT 177.425 105.320 177.700 106.170 ;
        RECT 177.420 105.150 177.700 105.320 ;
        RECT 177.425 105.010 177.700 105.150 ;
        RECT 177.870 104.810 178.060 106.170 ;
        RECT 178.240 105.805 178.750 106.340 ;
        RECT 178.970 105.530 179.215 106.135 ;
        RECT 180.670 105.790 180.840 106.170 ;
        RECT 181.055 105.960 181.385 106.340 ;
        RECT 180.670 105.620 181.385 105.790 ;
        RECT 178.260 105.360 179.490 105.530 ;
        RECT 177.050 104.640 178.060 104.810 ;
        RECT 178.230 104.795 178.980 104.985 ;
        RECT 176.710 104.300 177.835 104.470 ;
        RECT 178.230 104.130 178.400 104.795 ;
        RECT 179.150 104.550 179.490 105.360 ;
        RECT 180.580 105.070 180.935 105.440 ;
        RECT 181.215 105.430 181.385 105.620 ;
        RECT 181.555 105.595 181.810 106.170 ;
        RECT 181.215 105.100 181.470 105.430 ;
        RECT 181.215 104.890 181.385 105.100 ;
        RECT 176.370 103.960 178.400 104.130 ;
        RECT 178.570 103.790 178.740 104.550 ;
        RECT 178.975 104.140 179.490 104.550 ;
        RECT 180.670 104.720 181.385 104.890 ;
        RECT 181.640 104.865 181.810 105.595 ;
        RECT 181.985 105.500 182.245 106.340 ;
        RECT 182.510 105.790 182.680 106.170 ;
        RECT 182.895 105.960 183.225 106.340 ;
        RECT 182.510 105.620 183.225 105.790 ;
        RECT 182.420 105.070 182.775 105.440 ;
        RECT 183.055 105.430 183.225 105.620 ;
        RECT 183.395 105.595 183.650 106.170 ;
        RECT 183.055 105.100 183.310 105.430 ;
        RECT 180.670 103.960 180.840 104.720 ;
        RECT 181.055 103.790 181.385 104.550 ;
        RECT 181.555 103.960 181.810 104.865 ;
        RECT 181.985 103.790 182.245 104.940 ;
        RECT 183.055 104.890 183.225 105.100 ;
        RECT 182.510 104.720 183.225 104.890 ;
        RECT 183.480 104.865 183.650 105.595 ;
        RECT 183.825 105.500 184.085 106.340 ;
        RECT 184.260 105.600 184.645 106.170 ;
        RECT 184.815 105.880 185.140 106.340 ;
        RECT 185.660 105.710 185.940 106.170 ;
        RECT 182.510 103.960 182.680 104.720 ;
        RECT 182.895 103.790 183.225 104.550 ;
        RECT 183.395 103.960 183.650 104.865 ;
        RECT 183.825 103.790 184.085 104.940 ;
        RECT 184.260 104.930 184.540 105.600 ;
        RECT 184.815 105.540 185.940 105.710 ;
        RECT 184.815 105.430 185.265 105.540 ;
        RECT 184.710 105.100 185.265 105.430 ;
        RECT 186.130 105.370 186.530 106.170 ;
        RECT 186.930 105.880 187.200 106.340 ;
        RECT 187.370 105.710 187.655 106.170 ;
        RECT 184.260 103.960 184.645 104.930 ;
        RECT 184.815 104.640 185.265 105.100 ;
        RECT 185.435 104.810 186.530 105.370 ;
        RECT 184.815 104.420 185.940 104.640 ;
        RECT 184.815 103.790 185.140 104.250 ;
        RECT 185.660 103.960 185.940 104.420 ;
        RECT 186.130 103.960 186.530 104.810 ;
        RECT 186.700 105.540 187.655 105.710 ;
        RECT 187.940 105.615 188.230 106.340 ;
        RECT 188.405 105.790 188.660 106.080 ;
        RECT 188.830 105.960 189.160 106.340 ;
        RECT 188.405 105.620 189.155 105.790 ;
        RECT 186.700 104.640 186.910 105.540 ;
        RECT 187.080 104.810 187.770 105.370 ;
        RECT 186.700 104.420 187.655 104.640 ;
        RECT 186.930 103.790 187.200 104.250 ;
        RECT 187.370 103.960 187.655 104.420 ;
        RECT 187.940 103.790 188.230 104.955 ;
        RECT 188.405 104.800 188.755 105.450 ;
        RECT 188.925 104.630 189.155 105.620 ;
        RECT 188.405 104.460 189.155 104.630 ;
        RECT 188.405 103.960 188.660 104.460 ;
        RECT 188.830 103.790 189.160 104.290 ;
        RECT 189.330 103.960 189.500 106.080 ;
        RECT 189.860 105.980 190.190 106.340 ;
        RECT 190.360 105.950 190.855 106.120 ;
        RECT 191.060 105.950 191.915 106.120 ;
        RECT 189.730 104.760 190.190 105.810 ;
        RECT 189.670 103.975 189.995 104.760 ;
        RECT 190.360 104.590 190.530 105.950 ;
        RECT 190.700 105.040 191.050 105.660 ;
        RECT 191.220 105.440 191.575 105.660 ;
        RECT 191.220 104.850 191.390 105.440 ;
        RECT 191.745 105.240 191.915 105.950 ;
        RECT 192.790 105.880 193.120 106.340 ;
        RECT 193.330 105.980 193.680 106.150 ;
        RECT 192.120 105.410 192.910 105.660 ;
        RECT 193.330 105.590 193.590 105.980 ;
        RECT 193.900 105.890 194.850 106.170 ;
        RECT 195.020 105.900 195.210 106.340 ;
        RECT 195.380 105.960 196.450 106.130 ;
        RECT 193.080 105.240 193.250 105.420 ;
        RECT 190.360 104.420 190.755 104.590 ;
        RECT 190.925 104.460 191.390 104.850 ;
        RECT 191.560 105.070 193.250 105.240 ;
        RECT 190.585 104.290 190.755 104.420 ;
        RECT 191.560 104.290 191.730 105.070 ;
        RECT 193.420 104.900 193.590 105.590 ;
        RECT 192.090 104.730 193.590 104.900 ;
        RECT 193.780 104.930 193.990 105.720 ;
        RECT 194.160 105.100 194.510 105.720 ;
        RECT 194.680 105.110 194.850 105.890 ;
        RECT 195.380 105.730 195.550 105.960 ;
        RECT 195.020 105.560 195.550 105.730 ;
        RECT 195.020 105.280 195.240 105.560 ;
        RECT 195.720 105.390 195.960 105.790 ;
        RECT 194.680 104.940 195.085 105.110 ;
        RECT 195.420 105.020 195.960 105.390 ;
        RECT 196.130 105.605 196.450 105.960 ;
        RECT 196.695 105.880 197.000 106.340 ;
        RECT 197.170 105.630 197.425 106.160 ;
        RECT 196.130 105.430 196.455 105.605 ;
        RECT 196.130 105.130 197.045 105.430 ;
        RECT 196.305 105.100 197.045 105.130 ;
        RECT 193.780 104.770 194.455 104.930 ;
        RECT 194.915 104.850 195.085 104.940 ;
        RECT 193.780 104.760 194.745 104.770 ;
        RECT 193.420 104.590 193.590 104.730 ;
        RECT 190.165 103.790 190.415 104.250 ;
        RECT 190.585 103.960 190.835 104.290 ;
        RECT 191.050 103.960 191.730 104.290 ;
        RECT 191.900 104.390 192.975 104.560 ;
        RECT 193.420 104.420 193.980 104.590 ;
        RECT 194.285 104.470 194.745 104.760 ;
        RECT 194.915 104.680 196.135 104.850 ;
        RECT 191.900 104.050 192.070 104.390 ;
        RECT 192.305 103.790 192.635 104.220 ;
        RECT 192.805 104.050 192.975 104.390 ;
        RECT 193.270 103.790 193.640 104.250 ;
        RECT 193.810 103.960 193.980 104.420 ;
        RECT 194.915 104.300 195.085 104.680 ;
        RECT 196.305 104.510 196.475 105.100 ;
        RECT 197.215 104.980 197.425 105.630 ;
        RECT 197.600 105.590 198.810 106.340 ;
        RECT 199.070 105.790 199.240 106.170 ;
        RECT 199.455 105.960 199.785 106.340 ;
        RECT 199.070 105.620 199.785 105.790 ;
        RECT 197.600 105.050 198.120 105.590 ;
        RECT 194.215 103.960 195.085 104.300 ;
        RECT 195.675 104.340 196.475 104.510 ;
        RECT 195.255 103.790 195.505 104.250 ;
        RECT 195.675 104.050 195.845 104.340 ;
        RECT 196.025 103.790 196.355 104.170 ;
        RECT 196.695 103.790 197.000 104.930 ;
        RECT 197.170 104.100 197.425 104.980 ;
        RECT 198.290 104.880 198.810 105.420 ;
        RECT 198.980 105.070 199.335 105.440 ;
        RECT 199.615 105.430 199.785 105.620 ;
        RECT 199.955 105.595 200.210 106.170 ;
        RECT 199.615 105.100 199.870 105.430 ;
        RECT 199.615 104.890 199.785 105.100 ;
        RECT 197.600 103.790 198.810 104.880 ;
        RECT 199.070 104.720 199.785 104.890 ;
        RECT 200.040 104.865 200.210 105.595 ;
        RECT 200.385 105.500 200.645 106.340 ;
        RECT 200.820 105.615 201.110 106.340 ;
        RECT 201.370 105.790 201.540 106.170 ;
        RECT 201.755 105.960 202.085 106.340 ;
        RECT 201.370 105.620 202.085 105.790 ;
        RECT 201.280 105.070 201.635 105.440 ;
        RECT 201.915 105.430 202.085 105.620 ;
        RECT 202.255 105.595 202.510 106.170 ;
        RECT 201.915 105.100 202.170 105.430 ;
        RECT 199.070 103.960 199.240 104.720 ;
        RECT 199.455 103.790 199.785 104.550 ;
        RECT 199.955 103.960 200.210 104.865 ;
        RECT 200.385 103.790 200.645 104.940 ;
        RECT 200.820 103.790 201.110 104.955 ;
        RECT 201.915 104.890 202.085 105.100 ;
        RECT 201.370 104.720 202.085 104.890 ;
        RECT 202.340 104.865 202.510 105.595 ;
        RECT 202.685 105.500 202.945 106.340 ;
        RECT 203.210 105.790 203.380 106.170 ;
        RECT 203.595 105.960 203.925 106.340 ;
        RECT 203.210 105.620 203.925 105.790 ;
        RECT 203.120 105.070 203.475 105.440 ;
        RECT 203.755 105.430 203.925 105.620 ;
        RECT 204.095 105.595 204.350 106.170 ;
        RECT 203.755 105.100 204.010 105.430 ;
        RECT 201.370 103.960 201.540 104.720 ;
        RECT 201.755 103.790 202.085 104.550 ;
        RECT 202.255 103.960 202.510 104.865 ;
        RECT 202.685 103.790 202.945 104.940 ;
        RECT 203.755 104.890 203.925 105.100 ;
        RECT 203.210 104.720 203.925 104.890 ;
        RECT 204.180 104.865 204.350 105.595 ;
        RECT 204.525 105.500 204.785 106.340 ;
        RECT 204.965 105.500 205.225 106.340 ;
        RECT 205.400 105.595 205.655 106.170 ;
        RECT 205.825 105.960 206.155 106.340 ;
        RECT 206.370 105.790 206.540 106.170 ;
        RECT 205.825 105.620 206.540 105.790 ;
        RECT 203.210 103.960 203.380 104.720 ;
        RECT 203.595 103.790 203.925 104.550 ;
        RECT 204.095 103.960 204.350 104.865 ;
        RECT 204.525 103.790 204.785 104.940 ;
        RECT 204.965 103.790 205.225 104.940 ;
        RECT 205.400 104.865 205.570 105.595 ;
        RECT 205.825 105.430 205.995 105.620 ;
        RECT 206.805 105.600 207.060 106.170 ;
        RECT 207.230 105.940 207.560 106.340 ;
        RECT 207.985 105.805 208.515 106.170 ;
        RECT 207.985 105.770 208.160 105.805 ;
        RECT 207.230 105.600 208.160 105.770 ;
        RECT 205.740 105.100 205.995 105.430 ;
        RECT 205.825 104.890 205.995 105.100 ;
        RECT 206.275 105.070 206.630 105.440 ;
        RECT 206.805 104.930 206.975 105.600 ;
        RECT 207.230 105.430 207.400 105.600 ;
        RECT 207.145 105.100 207.400 105.430 ;
        RECT 207.625 105.100 207.820 105.430 ;
        RECT 205.400 103.960 205.655 104.865 ;
        RECT 205.825 104.720 206.540 104.890 ;
        RECT 205.825 103.790 206.155 104.550 ;
        RECT 206.370 103.960 206.540 104.720 ;
        RECT 206.805 103.960 207.140 104.930 ;
        RECT 207.310 103.790 207.480 104.930 ;
        RECT 207.650 104.130 207.820 105.100 ;
        RECT 207.990 104.470 208.160 105.600 ;
        RECT 208.330 104.810 208.500 105.610 ;
        RECT 208.705 105.320 208.980 106.170 ;
        RECT 208.700 105.150 208.980 105.320 ;
        RECT 208.705 105.010 208.980 105.150 ;
        RECT 209.150 104.810 209.340 106.170 ;
        RECT 209.520 105.805 210.030 106.340 ;
        RECT 210.250 105.530 210.495 106.135 ;
        RECT 209.540 105.360 210.770 105.530 ;
        RECT 211.865 105.500 212.125 106.340 ;
        RECT 212.300 105.595 212.555 106.170 ;
        RECT 212.725 105.960 213.055 106.340 ;
        RECT 213.270 105.790 213.440 106.170 ;
        RECT 212.725 105.620 213.440 105.790 ;
        RECT 208.330 104.640 209.340 104.810 ;
        RECT 209.510 104.795 210.260 104.985 ;
        RECT 207.990 104.300 209.115 104.470 ;
        RECT 209.510 104.130 209.680 104.795 ;
        RECT 210.430 104.550 210.770 105.360 ;
        RECT 207.650 103.960 209.680 104.130 ;
        RECT 209.850 103.790 210.020 104.550 ;
        RECT 210.255 104.140 210.770 104.550 ;
        RECT 211.865 103.790 212.125 104.940 ;
        RECT 212.300 104.865 212.470 105.595 ;
        RECT 212.725 105.430 212.895 105.620 ;
        RECT 213.700 105.615 213.990 106.340 ;
        RECT 214.165 105.500 214.425 106.340 ;
        RECT 214.600 105.595 214.855 106.170 ;
        RECT 215.025 105.960 215.355 106.340 ;
        RECT 215.570 105.790 215.740 106.170 ;
        RECT 215.025 105.620 215.740 105.790 ;
        RECT 212.640 105.100 212.895 105.430 ;
        RECT 212.725 104.890 212.895 105.100 ;
        RECT 213.175 105.070 213.530 105.440 ;
        RECT 212.300 103.960 212.555 104.865 ;
        RECT 212.725 104.720 213.440 104.890 ;
        RECT 212.725 103.790 213.055 104.550 ;
        RECT 213.270 103.960 213.440 104.720 ;
        RECT 213.700 103.790 213.990 104.955 ;
        RECT 214.165 103.790 214.425 104.940 ;
        RECT 214.600 104.865 214.770 105.595 ;
        RECT 215.025 105.430 215.195 105.620 ;
        RECT 216.005 105.500 216.265 106.340 ;
        RECT 216.440 105.595 216.695 106.170 ;
        RECT 216.865 105.960 217.195 106.340 ;
        RECT 217.410 105.790 217.580 106.170 ;
        RECT 216.865 105.620 217.580 105.790 ;
        RECT 217.930 105.790 218.100 106.170 ;
        RECT 218.315 105.960 218.645 106.340 ;
        RECT 217.930 105.620 218.645 105.790 ;
        RECT 214.940 105.100 215.195 105.430 ;
        RECT 215.025 104.890 215.195 105.100 ;
        RECT 215.475 105.070 215.830 105.440 ;
        RECT 214.600 103.960 214.855 104.865 ;
        RECT 215.025 104.720 215.740 104.890 ;
        RECT 215.025 103.790 215.355 104.550 ;
        RECT 215.570 103.960 215.740 104.720 ;
        RECT 216.005 103.790 216.265 104.940 ;
        RECT 216.440 104.865 216.610 105.595 ;
        RECT 216.865 105.430 217.035 105.620 ;
        RECT 216.780 105.100 217.035 105.430 ;
        RECT 216.865 104.890 217.035 105.100 ;
        RECT 217.315 105.070 217.670 105.440 ;
        RECT 217.840 105.070 218.195 105.440 ;
        RECT 218.475 105.430 218.645 105.620 ;
        RECT 218.815 105.595 219.070 106.170 ;
        RECT 218.475 105.100 218.730 105.430 ;
        RECT 218.475 104.890 218.645 105.100 ;
        RECT 216.440 103.960 216.695 104.865 ;
        RECT 216.865 104.720 217.580 104.890 ;
        RECT 216.865 103.790 217.195 104.550 ;
        RECT 217.410 103.960 217.580 104.720 ;
        RECT 217.930 104.720 218.645 104.890 ;
        RECT 218.900 104.865 219.070 105.595 ;
        RECT 219.245 105.500 219.505 106.340 ;
        RECT 219.685 105.600 219.940 106.170 ;
        RECT 220.110 105.940 220.440 106.340 ;
        RECT 220.865 105.805 221.395 106.170 ;
        RECT 220.865 105.770 221.040 105.805 ;
        RECT 220.110 105.600 221.040 105.770 ;
        RECT 221.585 105.660 221.860 106.170 ;
        RECT 217.930 103.960 218.100 104.720 ;
        RECT 218.315 103.790 218.645 104.550 ;
        RECT 218.815 103.960 219.070 104.865 ;
        RECT 219.245 103.790 219.505 104.940 ;
        RECT 219.685 104.930 219.855 105.600 ;
        RECT 220.110 105.430 220.280 105.600 ;
        RECT 220.025 105.100 220.280 105.430 ;
        RECT 220.505 105.100 220.700 105.430 ;
        RECT 219.685 103.960 220.020 104.930 ;
        RECT 220.190 103.790 220.360 104.930 ;
        RECT 220.530 104.130 220.700 105.100 ;
        RECT 220.870 104.470 221.040 105.600 ;
        RECT 221.210 104.810 221.380 105.610 ;
        RECT 221.580 105.490 221.860 105.660 ;
        RECT 221.585 105.010 221.860 105.490 ;
        RECT 222.030 104.810 222.220 106.170 ;
        RECT 222.400 105.805 222.910 106.340 ;
        RECT 223.130 105.530 223.375 106.135 ;
        RECT 222.420 105.360 223.650 105.530 ;
        RECT 224.745 105.500 225.005 106.340 ;
        RECT 225.180 105.595 225.435 106.170 ;
        RECT 225.605 105.960 225.935 106.340 ;
        RECT 226.150 105.790 226.320 106.170 ;
        RECT 225.605 105.620 226.320 105.790 ;
        RECT 221.210 104.640 222.220 104.810 ;
        RECT 222.390 104.795 223.140 104.985 ;
        RECT 220.870 104.300 221.995 104.470 ;
        RECT 222.390 104.130 222.560 104.795 ;
        RECT 223.310 104.550 223.650 105.360 ;
        RECT 220.530 103.960 222.560 104.130 ;
        RECT 222.730 103.790 222.900 104.550 ;
        RECT 223.135 104.140 223.650 104.550 ;
        RECT 224.745 103.790 225.005 104.940 ;
        RECT 225.180 104.865 225.350 105.595 ;
        RECT 225.605 105.430 225.775 105.620 ;
        RECT 226.580 105.615 226.870 106.340 ;
        RECT 227.040 105.600 227.425 106.170 ;
        RECT 227.595 105.880 227.920 106.340 ;
        RECT 228.440 105.710 228.720 106.170 ;
        RECT 225.520 105.100 225.775 105.430 ;
        RECT 225.605 104.890 225.775 105.100 ;
        RECT 226.055 105.070 226.410 105.440 ;
        RECT 225.180 103.960 225.435 104.865 ;
        RECT 225.605 104.720 226.320 104.890 ;
        RECT 225.605 103.790 225.935 104.550 ;
        RECT 226.150 103.960 226.320 104.720 ;
        RECT 226.580 103.790 226.870 104.955 ;
        RECT 227.040 104.930 227.320 105.600 ;
        RECT 227.595 105.540 228.720 105.710 ;
        RECT 227.595 105.430 228.045 105.540 ;
        RECT 227.490 105.100 228.045 105.430 ;
        RECT 228.910 105.370 229.310 106.170 ;
        RECT 229.710 105.880 229.980 106.340 ;
        RECT 230.150 105.710 230.435 106.170 ;
        RECT 227.040 103.960 227.425 104.930 ;
        RECT 227.595 104.640 228.045 105.100 ;
        RECT 228.215 104.810 229.310 105.370 ;
        RECT 227.595 104.420 228.720 104.640 ;
        RECT 227.595 103.790 227.920 104.250 ;
        RECT 228.440 103.960 228.720 104.420 ;
        RECT 228.910 103.960 229.310 104.810 ;
        RECT 229.480 105.540 230.435 105.710 ;
        RECT 229.480 104.640 229.690 105.540 ;
        RECT 231.185 105.500 231.445 106.340 ;
        RECT 231.620 105.595 231.875 106.170 ;
        RECT 232.045 105.960 232.375 106.340 ;
        RECT 232.590 105.790 232.760 106.170 ;
        RECT 232.045 105.620 232.760 105.790 ;
        RECT 229.860 104.810 230.550 105.370 ;
        RECT 229.480 104.420 230.435 104.640 ;
        RECT 229.710 103.790 229.980 104.250 ;
        RECT 230.150 103.960 230.435 104.420 ;
        RECT 231.185 103.790 231.445 104.940 ;
        RECT 231.620 104.865 231.790 105.595 ;
        RECT 232.045 105.430 232.215 105.620 ;
        RECT 233.485 105.500 233.745 106.340 ;
        RECT 233.920 105.595 234.175 106.170 ;
        RECT 234.345 105.960 234.675 106.340 ;
        RECT 234.890 105.790 235.060 106.170 ;
        RECT 234.345 105.620 235.060 105.790 ;
        RECT 235.870 105.790 236.040 106.170 ;
        RECT 236.255 105.960 236.585 106.340 ;
        RECT 235.870 105.620 236.585 105.790 ;
        RECT 231.960 105.100 232.215 105.430 ;
        RECT 232.045 104.890 232.215 105.100 ;
        RECT 232.495 105.070 232.850 105.440 ;
        RECT 231.620 103.960 231.875 104.865 ;
        RECT 232.045 104.720 232.760 104.890 ;
        RECT 232.045 103.790 232.375 104.550 ;
        RECT 232.590 103.960 232.760 104.720 ;
        RECT 233.485 103.790 233.745 104.940 ;
        RECT 233.920 104.865 234.090 105.595 ;
        RECT 234.345 105.430 234.515 105.620 ;
        RECT 234.260 105.100 234.515 105.430 ;
        RECT 234.345 104.890 234.515 105.100 ;
        RECT 234.795 105.070 235.150 105.440 ;
        RECT 235.780 105.070 236.135 105.440 ;
        RECT 236.415 105.430 236.585 105.620 ;
        RECT 236.755 105.595 237.010 106.170 ;
        RECT 236.415 105.100 236.670 105.430 ;
        RECT 236.415 104.890 236.585 105.100 ;
        RECT 233.920 103.960 234.175 104.865 ;
        RECT 234.345 104.720 235.060 104.890 ;
        RECT 234.345 103.790 234.675 104.550 ;
        RECT 234.890 103.960 235.060 104.720 ;
        RECT 235.870 104.720 236.585 104.890 ;
        RECT 236.840 104.865 237.010 105.595 ;
        RECT 237.185 105.500 237.445 106.340 ;
        RECT 237.625 105.500 237.885 106.340 ;
        RECT 238.060 105.595 238.315 106.170 ;
        RECT 238.485 105.960 238.815 106.340 ;
        RECT 239.030 105.790 239.200 106.170 ;
        RECT 238.485 105.620 239.200 105.790 ;
        RECT 235.870 103.960 236.040 104.720 ;
        RECT 236.255 103.790 236.585 104.550 ;
        RECT 236.755 103.960 237.010 104.865 ;
        RECT 237.185 103.790 237.445 104.940 ;
        RECT 237.625 103.790 237.885 104.940 ;
        RECT 238.060 104.865 238.230 105.595 ;
        RECT 238.485 105.430 238.655 105.620 ;
        RECT 239.460 105.615 239.750 106.340 ;
        RECT 239.925 105.600 240.180 106.170 ;
        RECT 240.350 105.940 240.680 106.340 ;
        RECT 241.105 105.805 241.635 106.170 ;
        RECT 241.105 105.770 241.280 105.805 ;
        RECT 240.350 105.600 241.280 105.770 ;
        RECT 238.400 105.100 238.655 105.430 ;
        RECT 238.485 104.890 238.655 105.100 ;
        RECT 238.935 105.070 239.290 105.440 ;
        RECT 238.060 103.960 238.315 104.865 ;
        RECT 238.485 104.720 239.200 104.890 ;
        RECT 238.485 103.790 238.815 104.550 ;
        RECT 239.030 103.960 239.200 104.720 ;
        RECT 239.460 103.790 239.750 104.955 ;
        RECT 239.925 104.930 240.095 105.600 ;
        RECT 240.350 105.430 240.520 105.600 ;
        RECT 240.265 105.100 240.520 105.430 ;
        RECT 240.745 105.100 240.940 105.430 ;
        RECT 239.925 103.960 240.260 104.930 ;
        RECT 240.430 103.790 240.600 104.930 ;
        RECT 240.770 104.130 240.940 105.100 ;
        RECT 241.110 104.470 241.280 105.600 ;
        RECT 241.450 104.810 241.620 105.610 ;
        RECT 241.825 105.320 242.100 106.170 ;
        RECT 241.820 105.150 242.100 105.320 ;
        RECT 241.825 105.010 242.100 105.150 ;
        RECT 242.270 104.810 242.460 106.170 ;
        RECT 242.640 105.805 243.150 106.340 ;
        RECT 243.370 105.530 243.615 106.135 ;
        RECT 244.060 105.600 244.445 106.170 ;
        RECT 244.615 105.880 244.940 106.340 ;
        RECT 245.460 105.710 245.740 106.170 ;
        RECT 242.660 105.360 243.890 105.530 ;
        RECT 241.450 104.640 242.460 104.810 ;
        RECT 242.630 104.795 243.380 104.985 ;
        RECT 241.110 104.300 242.235 104.470 ;
        RECT 242.630 104.130 242.800 104.795 ;
        RECT 243.550 104.550 243.890 105.360 ;
        RECT 240.770 103.960 242.800 104.130 ;
        RECT 242.970 103.790 243.140 104.550 ;
        RECT 243.375 104.140 243.890 104.550 ;
        RECT 244.060 104.930 244.340 105.600 ;
        RECT 244.615 105.540 245.740 105.710 ;
        RECT 244.615 105.430 245.065 105.540 ;
        RECT 244.510 105.100 245.065 105.430 ;
        RECT 245.930 105.370 246.330 106.170 ;
        RECT 246.730 105.880 247.000 106.340 ;
        RECT 247.170 105.710 247.455 106.170 ;
        RECT 244.060 103.960 244.445 104.930 ;
        RECT 244.615 104.640 245.065 105.100 ;
        RECT 245.235 104.810 246.330 105.370 ;
        RECT 244.615 104.420 245.740 104.640 ;
        RECT 244.615 103.790 244.940 104.250 ;
        RECT 245.460 103.960 245.740 104.420 ;
        RECT 245.930 103.960 246.330 104.810 ;
        RECT 246.500 105.540 247.455 105.710 ;
        RECT 247.740 105.600 248.125 106.170 ;
        RECT 248.295 105.880 248.620 106.340 ;
        RECT 249.140 105.710 249.420 106.170 ;
        RECT 246.500 104.640 246.710 105.540 ;
        RECT 246.880 104.810 247.570 105.370 ;
        RECT 247.740 104.930 248.020 105.600 ;
        RECT 248.295 105.540 249.420 105.710 ;
        RECT 248.295 105.430 248.745 105.540 ;
        RECT 248.190 105.100 248.745 105.430 ;
        RECT 249.610 105.370 250.010 106.170 ;
        RECT 250.410 105.880 250.680 106.340 ;
        RECT 250.850 105.710 251.135 106.170 ;
        RECT 246.500 104.420 247.455 104.640 ;
        RECT 246.730 103.790 247.000 104.250 ;
        RECT 247.170 103.960 247.455 104.420 ;
        RECT 247.740 103.960 248.125 104.930 ;
        RECT 248.295 104.640 248.745 105.100 ;
        RECT 248.915 104.810 250.010 105.370 ;
        RECT 248.295 104.420 249.420 104.640 ;
        RECT 248.295 103.790 248.620 104.250 ;
        RECT 249.140 103.960 249.420 104.420 ;
        RECT 249.610 103.960 250.010 104.810 ;
        RECT 250.180 105.540 251.135 105.710 ;
        RECT 252.340 105.615 252.630 106.340 ;
        RECT 252.915 105.710 253.200 106.170 ;
        RECT 253.370 105.880 253.640 106.340 ;
        RECT 252.915 105.540 253.870 105.710 ;
        RECT 250.180 104.640 250.390 105.540 ;
        RECT 250.560 104.810 251.250 105.370 ;
        RECT 250.180 104.420 251.135 104.640 ;
        RECT 250.410 103.790 250.680 104.250 ;
        RECT 250.850 103.960 251.135 104.420 ;
        RECT 252.340 103.790 252.630 104.955 ;
        RECT 252.800 104.810 253.490 105.370 ;
        RECT 253.660 104.640 253.870 105.540 ;
        RECT 252.915 104.420 253.870 104.640 ;
        RECT 254.040 105.370 254.440 106.170 ;
        RECT 254.630 105.710 254.910 106.170 ;
        RECT 255.430 105.880 255.755 106.340 ;
        RECT 254.630 105.540 255.755 105.710 ;
        RECT 255.925 105.600 256.310 106.170 ;
        RECT 255.305 105.430 255.755 105.540 ;
        RECT 254.040 104.810 255.135 105.370 ;
        RECT 255.305 105.100 255.860 105.430 ;
        RECT 252.915 103.960 253.200 104.420 ;
        RECT 253.370 103.790 253.640 104.250 ;
        RECT 254.040 103.960 254.440 104.810 ;
        RECT 255.305 104.640 255.755 105.100 ;
        RECT 256.030 104.930 256.310 105.600 ;
        RECT 254.630 104.420 255.755 104.640 ;
        RECT 254.630 103.960 254.910 104.420 ;
        RECT 255.430 103.790 255.755 104.250 ;
        RECT 255.925 103.960 256.310 104.930 ;
        RECT 257.405 105.600 257.660 106.170 ;
        RECT 257.830 105.940 258.160 106.340 ;
        RECT 258.585 105.805 259.115 106.170 ;
        RECT 258.585 105.770 258.760 105.805 ;
        RECT 257.830 105.600 258.760 105.770 ;
        RECT 257.405 104.930 257.575 105.600 ;
        RECT 257.830 105.430 258.000 105.600 ;
        RECT 257.745 105.100 258.000 105.430 ;
        RECT 258.225 105.100 258.420 105.430 ;
        RECT 257.405 103.960 257.740 104.930 ;
        RECT 257.910 103.790 258.080 104.930 ;
        RECT 258.250 104.130 258.420 105.100 ;
        RECT 258.590 104.470 258.760 105.600 ;
        RECT 258.930 104.810 259.100 105.610 ;
        RECT 259.305 105.320 259.580 106.170 ;
        RECT 259.300 105.150 259.580 105.320 ;
        RECT 259.305 105.010 259.580 105.150 ;
        RECT 259.750 104.810 259.940 106.170 ;
        RECT 260.120 105.805 260.630 106.340 ;
        RECT 260.850 105.530 261.095 106.135 ;
        RECT 261.630 105.790 261.800 106.170 ;
        RECT 262.015 105.960 262.345 106.340 ;
        RECT 261.630 105.620 262.345 105.790 ;
        RECT 260.140 105.360 261.370 105.530 ;
        RECT 258.930 104.640 259.940 104.810 ;
        RECT 260.110 104.795 260.860 104.985 ;
        RECT 258.590 104.300 259.715 104.470 ;
        RECT 260.110 104.130 260.280 104.795 ;
        RECT 261.030 104.550 261.370 105.360 ;
        RECT 261.540 105.070 261.895 105.440 ;
        RECT 262.175 105.430 262.345 105.620 ;
        RECT 262.515 105.595 262.770 106.170 ;
        RECT 262.175 105.100 262.430 105.430 ;
        RECT 262.175 104.890 262.345 105.100 ;
        RECT 258.250 103.960 260.280 104.130 ;
        RECT 260.450 103.790 260.620 104.550 ;
        RECT 260.855 104.140 261.370 104.550 ;
        RECT 261.630 104.720 262.345 104.890 ;
        RECT 262.600 104.865 262.770 105.595 ;
        RECT 262.945 105.500 263.205 106.340 ;
        RECT 263.470 105.790 263.640 106.170 ;
        RECT 263.855 105.960 264.185 106.340 ;
        RECT 263.470 105.620 264.185 105.790 ;
        RECT 263.380 105.070 263.735 105.440 ;
        RECT 264.015 105.430 264.185 105.620 ;
        RECT 264.355 105.595 264.610 106.170 ;
        RECT 264.015 105.100 264.270 105.430 ;
        RECT 261.630 103.960 261.800 104.720 ;
        RECT 262.015 103.790 262.345 104.550 ;
        RECT 262.515 103.960 262.770 104.865 ;
        RECT 262.945 103.790 263.205 104.940 ;
        RECT 264.015 104.890 264.185 105.100 ;
        RECT 263.470 104.720 264.185 104.890 ;
        RECT 264.440 104.865 264.610 105.595 ;
        RECT 264.785 105.500 265.045 106.340 ;
        RECT 265.220 105.615 265.510 106.340 ;
        RECT 265.685 105.500 265.945 106.340 ;
        RECT 266.120 105.595 266.375 106.170 ;
        RECT 266.545 105.960 266.875 106.340 ;
        RECT 267.090 105.790 267.260 106.170 ;
        RECT 266.545 105.620 267.260 105.790 ;
        RECT 263.470 103.960 263.640 104.720 ;
        RECT 263.855 103.790 264.185 104.550 ;
        RECT 264.355 103.960 264.610 104.865 ;
        RECT 264.785 103.790 265.045 104.940 ;
        RECT 265.220 103.790 265.510 104.955 ;
        RECT 265.685 103.790 265.945 104.940 ;
        RECT 266.120 104.865 266.290 105.595 ;
        RECT 266.545 105.430 266.715 105.620 ;
        RECT 267.525 105.500 267.785 106.340 ;
        RECT 267.960 105.595 268.215 106.170 ;
        RECT 268.385 105.960 268.715 106.340 ;
        RECT 268.930 105.790 269.100 106.170 ;
        RECT 268.385 105.620 269.100 105.790 ;
        RECT 266.460 105.100 266.715 105.430 ;
        RECT 266.545 104.890 266.715 105.100 ;
        RECT 266.995 105.070 267.350 105.440 ;
        RECT 266.120 103.960 266.375 104.865 ;
        RECT 266.545 104.720 267.260 104.890 ;
        RECT 266.545 103.790 266.875 104.550 ;
        RECT 267.090 103.960 267.260 104.720 ;
        RECT 267.525 103.790 267.785 104.940 ;
        RECT 267.960 104.865 268.130 105.595 ;
        RECT 268.385 105.430 268.555 105.620 ;
        RECT 269.365 105.500 269.625 106.340 ;
        RECT 269.800 105.595 270.055 106.170 ;
        RECT 270.225 105.960 270.555 106.340 ;
        RECT 270.770 105.790 270.940 106.170 ;
        RECT 270.225 105.620 270.940 105.790 ;
        RECT 268.300 105.100 268.555 105.430 ;
        RECT 268.385 104.890 268.555 105.100 ;
        RECT 268.835 105.070 269.190 105.440 ;
        RECT 267.960 103.960 268.215 104.865 ;
        RECT 268.385 104.720 269.100 104.890 ;
        RECT 268.385 103.790 268.715 104.550 ;
        RECT 268.930 103.960 269.100 104.720 ;
        RECT 269.365 103.790 269.625 104.940 ;
        RECT 269.800 104.865 269.970 105.595 ;
        RECT 270.225 105.430 270.395 105.620 ;
        RECT 271.200 105.590 272.410 106.340 ;
        RECT 272.580 105.600 272.965 106.170 ;
        RECT 273.135 105.880 273.460 106.340 ;
        RECT 273.980 105.710 274.260 106.170 ;
        RECT 270.140 105.100 270.395 105.430 ;
        RECT 270.225 104.890 270.395 105.100 ;
        RECT 270.675 105.070 271.030 105.440 ;
        RECT 271.200 105.050 271.720 105.590 ;
        RECT 269.800 103.960 270.055 104.865 ;
        RECT 270.225 104.720 270.940 104.890 ;
        RECT 271.890 104.880 272.410 105.420 ;
        RECT 270.225 103.790 270.555 104.550 ;
        RECT 270.770 103.960 270.940 104.720 ;
        RECT 271.200 103.790 272.410 104.880 ;
        RECT 272.580 104.930 272.860 105.600 ;
        RECT 273.135 105.540 274.260 105.710 ;
        RECT 273.135 105.430 273.585 105.540 ;
        RECT 273.030 105.100 273.585 105.430 ;
        RECT 274.450 105.370 274.850 106.170 ;
        RECT 275.250 105.880 275.520 106.340 ;
        RECT 275.690 105.710 275.975 106.170 ;
        RECT 272.580 103.960 272.965 104.930 ;
        RECT 273.135 104.640 273.585 105.100 ;
        RECT 273.755 104.810 274.850 105.370 ;
        RECT 273.135 104.420 274.260 104.640 ;
        RECT 273.135 103.790 273.460 104.250 ;
        RECT 273.980 103.960 274.260 104.420 ;
        RECT 274.450 103.960 274.850 104.810 ;
        RECT 275.020 105.540 275.975 105.710 ;
        RECT 275.020 104.640 275.230 105.540 ;
        RECT 276.265 105.500 276.525 106.340 ;
        RECT 276.700 105.595 276.955 106.170 ;
        RECT 277.125 105.960 277.455 106.340 ;
        RECT 277.670 105.790 277.840 106.170 ;
        RECT 277.125 105.620 277.840 105.790 ;
        RECT 275.400 104.810 276.090 105.370 ;
        RECT 275.020 104.420 275.975 104.640 ;
        RECT 275.250 103.790 275.520 104.250 ;
        RECT 275.690 103.960 275.975 104.420 ;
        RECT 276.265 103.790 276.525 104.940 ;
        RECT 276.700 104.865 276.870 105.595 ;
        RECT 277.125 105.430 277.295 105.620 ;
        RECT 278.100 105.615 278.390 106.340 ;
        RECT 278.565 105.630 278.820 106.160 ;
        RECT 278.990 105.880 279.295 106.340 ;
        RECT 279.540 105.960 280.610 106.130 ;
        RECT 277.040 105.100 277.295 105.430 ;
        RECT 277.125 104.890 277.295 105.100 ;
        RECT 277.575 105.070 277.930 105.440 ;
        RECT 278.565 104.980 278.775 105.630 ;
        RECT 279.540 105.605 279.860 105.960 ;
        RECT 279.535 105.430 279.860 105.605 ;
        RECT 278.945 105.130 279.860 105.430 ;
        RECT 280.030 105.390 280.270 105.790 ;
        RECT 280.440 105.730 280.610 105.960 ;
        RECT 280.780 105.900 280.970 106.340 ;
        RECT 281.140 105.890 282.090 106.170 ;
        RECT 282.310 105.980 282.660 106.150 ;
        RECT 280.440 105.560 280.970 105.730 ;
        RECT 278.945 105.100 279.685 105.130 ;
        RECT 276.700 103.960 276.955 104.865 ;
        RECT 277.125 104.720 277.840 104.890 ;
        RECT 277.125 103.790 277.455 104.550 ;
        RECT 277.670 103.960 277.840 104.720 ;
        RECT 278.100 103.790 278.390 104.955 ;
        RECT 278.565 104.100 278.820 104.980 ;
        RECT 278.990 103.790 279.295 104.930 ;
        RECT 279.515 104.510 279.685 105.100 ;
        RECT 280.030 105.020 280.570 105.390 ;
        RECT 280.750 105.280 280.970 105.560 ;
        RECT 281.140 105.110 281.310 105.890 ;
        RECT 280.905 104.940 281.310 105.110 ;
        RECT 281.480 105.100 281.830 105.720 ;
        RECT 280.905 104.850 281.075 104.940 ;
        RECT 282.000 104.930 282.210 105.720 ;
        RECT 279.855 104.680 281.075 104.850 ;
        RECT 281.535 104.770 282.210 104.930 ;
        RECT 279.515 104.340 280.315 104.510 ;
        RECT 279.635 103.790 279.965 104.170 ;
        RECT 280.145 104.050 280.315 104.340 ;
        RECT 280.905 104.300 281.075 104.680 ;
        RECT 281.245 104.760 282.210 104.770 ;
        RECT 282.400 105.590 282.660 105.980 ;
        RECT 282.870 105.880 283.200 106.340 ;
        RECT 284.075 105.950 284.930 106.120 ;
        RECT 285.135 105.950 285.630 106.120 ;
        RECT 285.800 105.980 286.130 106.340 ;
        RECT 282.400 104.900 282.570 105.590 ;
        RECT 282.740 105.240 282.910 105.420 ;
        RECT 283.080 105.410 283.870 105.660 ;
        RECT 284.075 105.240 284.245 105.950 ;
        RECT 284.415 105.440 284.770 105.660 ;
        RECT 282.740 105.070 284.430 105.240 ;
        RECT 281.245 104.470 281.705 104.760 ;
        RECT 282.400 104.730 283.900 104.900 ;
        RECT 282.400 104.590 282.570 104.730 ;
        RECT 282.010 104.420 282.570 104.590 ;
        RECT 280.485 103.790 280.735 104.250 ;
        RECT 280.905 103.960 281.775 104.300 ;
        RECT 282.010 103.960 282.180 104.420 ;
        RECT 283.015 104.390 284.090 104.560 ;
        RECT 282.350 103.790 282.720 104.250 ;
        RECT 283.015 104.050 283.185 104.390 ;
        RECT 283.355 103.790 283.685 104.220 ;
        RECT 283.920 104.050 284.090 104.390 ;
        RECT 284.260 104.290 284.430 105.070 ;
        RECT 284.600 104.850 284.770 105.440 ;
        RECT 284.940 105.040 285.290 105.660 ;
        RECT 284.600 104.460 285.065 104.850 ;
        RECT 285.460 104.590 285.630 105.950 ;
        RECT 285.800 104.760 286.260 105.810 ;
        RECT 285.235 104.420 285.630 104.590 ;
        RECT 285.235 104.290 285.405 104.420 ;
        RECT 284.260 103.960 284.940 104.290 ;
        RECT 285.155 103.960 285.405 104.290 ;
        RECT 285.575 103.790 285.825 104.250 ;
        RECT 285.995 103.975 286.320 104.760 ;
        RECT 286.490 103.960 286.660 106.080 ;
        RECT 286.830 105.960 287.160 106.340 ;
        RECT 287.330 105.790 287.585 106.080 ;
        RECT 286.835 105.620 287.585 105.790 ;
        RECT 286.835 104.630 287.065 105.620 ;
        RECT 287.765 105.500 288.025 106.340 ;
        RECT 288.200 105.595 288.455 106.170 ;
        RECT 288.625 105.960 288.955 106.340 ;
        RECT 289.170 105.790 289.340 106.170 ;
        RECT 288.625 105.620 289.340 105.790 ;
        RECT 287.235 104.800 287.585 105.450 ;
        RECT 286.835 104.460 287.585 104.630 ;
        RECT 286.830 103.790 287.160 104.290 ;
        RECT 287.330 103.960 287.585 104.460 ;
        RECT 287.765 103.790 288.025 104.940 ;
        RECT 288.200 104.865 288.370 105.595 ;
        RECT 288.625 105.430 288.795 105.620 ;
        RECT 289.600 105.590 290.810 106.340 ;
        RECT 290.980 105.615 291.270 106.340 ;
        RECT 288.540 105.100 288.795 105.430 ;
        RECT 288.625 104.890 288.795 105.100 ;
        RECT 289.075 105.070 289.430 105.440 ;
        RECT 289.600 105.050 290.120 105.590 ;
        RECT 291.445 105.500 291.705 106.340 ;
        RECT 291.880 105.595 292.135 106.170 ;
        RECT 292.305 105.960 292.635 106.340 ;
        RECT 292.850 105.790 293.020 106.170 ;
        RECT 292.305 105.620 293.020 105.790 ;
        RECT 288.200 103.960 288.455 104.865 ;
        RECT 288.625 104.720 289.340 104.890 ;
        RECT 290.290 104.880 290.810 105.420 ;
        RECT 288.625 103.790 288.955 104.550 ;
        RECT 289.170 103.960 289.340 104.720 ;
        RECT 289.600 103.790 290.810 104.880 ;
        RECT 290.980 103.790 291.270 104.955 ;
        RECT 291.445 103.790 291.705 104.940 ;
        RECT 291.880 104.865 292.050 105.595 ;
        RECT 292.305 105.430 292.475 105.620 ;
        RECT 293.280 105.590 294.490 106.340 ;
        RECT 294.665 105.790 294.920 106.080 ;
        RECT 295.090 105.960 295.420 106.340 ;
        RECT 294.665 105.620 295.415 105.790 ;
        RECT 292.220 105.100 292.475 105.430 ;
        RECT 292.305 104.890 292.475 105.100 ;
        RECT 292.755 105.070 293.110 105.440 ;
        RECT 293.280 105.050 293.800 105.590 ;
        RECT 291.880 103.960 292.135 104.865 ;
        RECT 292.305 104.720 293.020 104.890 ;
        RECT 293.970 104.880 294.490 105.420 ;
        RECT 292.305 103.790 292.635 104.550 ;
        RECT 292.850 103.960 293.020 104.720 ;
        RECT 293.280 103.790 294.490 104.880 ;
        RECT 294.665 104.800 295.015 105.450 ;
        RECT 295.185 104.630 295.415 105.620 ;
        RECT 294.665 104.460 295.415 104.630 ;
        RECT 294.665 103.960 294.920 104.460 ;
        RECT 295.090 103.790 295.420 104.290 ;
        RECT 295.590 103.960 295.760 106.080 ;
        RECT 296.120 105.980 296.450 106.340 ;
        RECT 296.620 105.950 297.115 106.120 ;
        RECT 297.320 105.950 298.175 106.120 ;
        RECT 295.990 104.760 296.450 105.810 ;
        RECT 295.930 103.975 296.255 104.760 ;
        RECT 296.620 104.590 296.790 105.950 ;
        RECT 296.960 105.040 297.310 105.660 ;
        RECT 297.480 105.440 297.835 105.660 ;
        RECT 297.480 104.850 297.650 105.440 ;
        RECT 298.005 105.240 298.175 105.950 ;
        RECT 299.050 105.880 299.380 106.340 ;
        RECT 299.590 105.980 299.940 106.150 ;
        RECT 298.380 105.410 299.170 105.660 ;
        RECT 299.590 105.590 299.850 105.980 ;
        RECT 300.160 105.890 301.110 106.170 ;
        RECT 301.280 105.900 301.470 106.340 ;
        RECT 301.640 105.960 302.710 106.130 ;
        RECT 299.340 105.240 299.510 105.420 ;
        RECT 296.620 104.420 297.015 104.590 ;
        RECT 297.185 104.460 297.650 104.850 ;
        RECT 297.820 105.070 299.510 105.240 ;
        RECT 296.845 104.290 297.015 104.420 ;
        RECT 297.820 104.290 297.990 105.070 ;
        RECT 299.680 104.900 299.850 105.590 ;
        RECT 298.350 104.730 299.850 104.900 ;
        RECT 300.040 104.930 300.250 105.720 ;
        RECT 300.420 105.100 300.770 105.720 ;
        RECT 300.940 105.110 301.110 105.890 ;
        RECT 301.640 105.730 301.810 105.960 ;
        RECT 301.280 105.560 301.810 105.730 ;
        RECT 301.280 105.280 301.500 105.560 ;
        RECT 301.980 105.390 302.220 105.790 ;
        RECT 300.940 104.940 301.345 105.110 ;
        RECT 301.680 105.020 302.220 105.390 ;
        RECT 302.390 105.605 302.710 105.960 ;
        RECT 302.955 105.880 303.260 106.340 ;
        RECT 303.430 105.630 303.685 106.160 ;
        RECT 302.390 105.430 302.715 105.605 ;
        RECT 302.390 105.130 303.305 105.430 ;
        RECT 302.565 105.100 303.305 105.130 ;
        RECT 300.040 104.770 300.715 104.930 ;
        RECT 301.175 104.850 301.345 104.940 ;
        RECT 300.040 104.760 301.005 104.770 ;
        RECT 299.680 104.590 299.850 104.730 ;
        RECT 296.425 103.790 296.675 104.250 ;
        RECT 296.845 103.960 297.095 104.290 ;
        RECT 297.310 103.960 297.990 104.290 ;
        RECT 298.160 104.390 299.235 104.560 ;
        RECT 299.680 104.420 300.240 104.590 ;
        RECT 300.545 104.470 301.005 104.760 ;
        RECT 301.175 104.680 302.395 104.850 ;
        RECT 298.160 104.050 298.330 104.390 ;
        RECT 298.565 103.790 298.895 104.220 ;
        RECT 299.065 104.050 299.235 104.390 ;
        RECT 299.530 103.790 299.900 104.250 ;
        RECT 300.070 103.960 300.240 104.420 ;
        RECT 301.175 104.300 301.345 104.680 ;
        RECT 302.565 104.510 302.735 105.100 ;
        RECT 303.475 104.980 303.685 105.630 ;
        RECT 303.860 105.615 304.150 106.340 ;
        RECT 304.325 105.500 304.585 106.340 ;
        RECT 304.760 105.595 305.015 106.170 ;
        RECT 305.185 105.960 305.515 106.340 ;
        RECT 305.730 105.790 305.900 106.170 ;
        RECT 305.185 105.620 305.900 105.790 ;
        RECT 307.170 105.790 307.340 106.170 ;
        RECT 307.555 105.960 307.885 106.340 ;
        RECT 307.170 105.620 307.885 105.790 ;
        RECT 300.475 103.960 301.345 104.300 ;
        RECT 301.935 104.340 302.735 104.510 ;
        RECT 301.515 103.790 301.765 104.250 ;
        RECT 301.935 104.050 302.105 104.340 ;
        RECT 302.285 103.790 302.615 104.170 ;
        RECT 302.955 103.790 303.260 104.930 ;
        RECT 303.430 104.100 303.685 104.980 ;
        RECT 303.860 103.790 304.150 104.955 ;
        RECT 304.325 103.790 304.585 104.940 ;
        RECT 304.760 104.865 304.930 105.595 ;
        RECT 305.185 105.430 305.355 105.620 ;
        RECT 305.100 105.100 305.355 105.430 ;
        RECT 305.185 104.890 305.355 105.100 ;
        RECT 305.635 105.070 305.990 105.440 ;
        RECT 307.080 105.070 307.435 105.440 ;
        RECT 307.715 105.430 307.885 105.620 ;
        RECT 308.055 105.595 308.310 106.170 ;
        RECT 307.715 105.100 307.970 105.430 ;
        RECT 307.715 104.890 307.885 105.100 ;
        RECT 304.760 103.960 305.015 104.865 ;
        RECT 305.185 104.720 305.900 104.890 ;
        RECT 305.185 103.790 305.515 104.550 ;
        RECT 305.730 103.960 305.900 104.720 ;
        RECT 307.170 104.720 307.885 104.890 ;
        RECT 308.140 104.865 308.310 105.595 ;
        RECT 308.485 105.500 308.745 106.340 ;
        RECT 309.840 105.590 311.050 106.340 ;
        RECT 307.170 103.960 307.340 104.720 ;
        RECT 307.555 103.790 307.885 104.550 ;
        RECT 308.055 103.960 308.310 104.865 ;
        RECT 308.485 103.790 308.745 104.940 ;
        RECT 309.840 104.880 310.360 105.420 ;
        RECT 310.530 105.050 311.050 105.590 ;
        RECT 309.840 103.790 311.050 104.880 ;
        RECT 162.095 103.620 311.135 103.790 ;
        RECT 162.180 102.530 163.390 103.620 ;
        RECT 162.180 101.820 162.700 102.360 ;
        RECT 162.870 101.990 163.390 102.530 ;
        RECT 164.025 102.470 164.285 103.620 ;
        RECT 164.460 102.545 164.715 103.450 ;
        RECT 164.885 102.860 165.215 103.620 ;
        RECT 165.430 102.690 165.600 103.450 ;
        RECT 165.865 102.950 166.120 103.450 ;
        RECT 166.290 103.120 166.620 103.620 ;
        RECT 165.865 102.780 166.615 102.950 ;
        RECT 162.180 101.070 163.390 101.820 ;
        RECT 164.025 101.070 164.285 101.910 ;
        RECT 164.460 101.815 164.630 102.545 ;
        RECT 164.885 102.520 165.600 102.690 ;
        RECT 164.885 102.310 165.055 102.520 ;
        RECT 164.800 101.980 165.055 102.310 ;
        RECT 164.460 101.240 164.715 101.815 ;
        RECT 164.885 101.790 165.055 101.980 ;
        RECT 165.335 101.970 165.690 102.340 ;
        RECT 165.865 101.960 166.215 102.610 ;
        RECT 166.385 101.790 166.615 102.780 ;
        RECT 164.885 101.620 165.600 101.790 ;
        RECT 164.885 101.070 165.215 101.450 ;
        RECT 165.430 101.240 165.600 101.620 ;
        RECT 165.865 101.620 166.615 101.790 ;
        RECT 165.865 101.330 166.120 101.620 ;
        RECT 166.290 101.070 166.620 101.450 ;
        RECT 166.790 101.330 166.960 103.450 ;
        RECT 167.130 102.650 167.455 103.435 ;
        RECT 167.625 103.160 167.875 103.620 ;
        RECT 168.045 103.120 168.295 103.450 ;
        RECT 168.510 103.120 169.190 103.450 ;
        RECT 168.045 102.990 168.215 103.120 ;
        RECT 167.820 102.820 168.215 102.990 ;
        RECT 167.190 101.600 167.650 102.650 ;
        RECT 167.820 101.460 167.990 102.820 ;
        RECT 168.385 102.560 168.850 102.950 ;
        RECT 168.160 101.750 168.510 102.370 ;
        RECT 168.680 101.970 168.850 102.560 ;
        RECT 169.020 102.340 169.190 103.120 ;
        RECT 169.360 103.020 169.530 103.360 ;
        RECT 169.765 103.190 170.095 103.620 ;
        RECT 170.265 103.020 170.435 103.360 ;
        RECT 170.730 103.160 171.100 103.620 ;
        RECT 169.360 102.850 170.435 103.020 ;
        RECT 171.270 102.990 171.440 103.450 ;
        RECT 171.675 103.110 172.545 103.450 ;
        RECT 172.715 103.160 172.965 103.620 ;
        RECT 170.880 102.820 171.440 102.990 ;
        RECT 170.880 102.680 171.050 102.820 ;
        RECT 169.550 102.510 171.050 102.680 ;
        RECT 171.745 102.650 172.205 102.940 ;
        RECT 169.020 102.170 170.710 102.340 ;
        RECT 168.680 101.750 169.035 101.970 ;
        RECT 169.205 101.460 169.375 102.170 ;
        RECT 169.580 101.750 170.370 102.000 ;
        RECT 170.540 101.990 170.710 102.170 ;
        RECT 170.880 101.820 171.050 102.510 ;
        RECT 167.320 101.070 167.650 101.430 ;
        RECT 167.820 101.290 168.315 101.460 ;
        RECT 168.520 101.290 169.375 101.460 ;
        RECT 170.250 101.070 170.580 101.530 ;
        RECT 170.790 101.430 171.050 101.820 ;
        RECT 171.240 102.640 172.205 102.650 ;
        RECT 172.375 102.730 172.545 103.110 ;
        RECT 173.135 103.070 173.305 103.360 ;
        RECT 173.485 103.240 173.815 103.620 ;
        RECT 173.135 102.900 173.935 103.070 ;
        RECT 171.240 102.480 171.915 102.640 ;
        RECT 172.375 102.560 173.595 102.730 ;
        RECT 171.240 101.690 171.450 102.480 ;
        RECT 172.375 102.470 172.545 102.560 ;
        RECT 171.620 101.690 171.970 102.310 ;
        RECT 172.140 102.300 172.545 102.470 ;
        RECT 172.140 101.520 172.310 102.300 ;
        RECT 172.480 101.850 172.700 102.130 ;
        RECT 172.880 102.020 173.420 102.390 ;
        RECT 173.765 102.310 173.935 102.900 ;
        RECT 174.155 102.480 174.460 103.620 ;
        RECT 174.630 102.430 174.885 103.310 ;
        RECT 175.060 102.455 175.350 103.620 ;
        RECT 175.525 102.950 175.780 103.450 ;
        RECT 175.950 103.120 176.280 103.620 ;
        RECT 175.525 102.780 176.275 102.950 ;
        RECT 173.765 102.280 174.505 102.310 ;
        RECT 172.480 101.680 173.010 101.850 ;
        RECT 170.790 101.260 171.140 101.430 ;
        RECT 171.360 101.240 172.310 101.520 ;
        RECT 172.480 101.070 172.670 101.510 ;
        RECT 172.840 101.450 173.010 101.680 ;
        RECT 173.180 101.620 173.420 102.020 ;
        RECT 173.590 101.980 174.505 102.280 ;
        RECT 173.590 101.805 173.915 101.980 ;
        RECT 173.590 101.450 173.910 101.805 ;
        RECT 174.675 101.780 174.885 102.430 ;
        RECT 175.525 101.960 175.875 102.610 ;
        RECT 172.840 101.280 173.910 101.450 ;
        RECT 174.155 101.070 174.460 101.530 ;
        RECT 174.630 101.250 174.885 101.780 ;
        RECT 175.060 101.070 175.350 101.795 ;
        RECT 176.045 101.790 176.275 102.780 ;
        RECT 175.525 101.620 176.275 101.790 ;
        RECT 175.525 101.330 175.780 101.620 ;
        RECT 175.950 101.070 176.280 101.450 ;
        RECT 176.450 101.330 176.620 103.450 ;
        RECT 176.790 102.650 177.115 103.435 ;
        RECT 177.285 103.160 177.535 103.620 ;
        RECT 177.705 103.120 177.955 103.450 ;
        RECT 178.170 103.120 178.850 103.450 ;
        RECT 177.705 102.990 177.875 103.120 ;
        RECT 177.480 102.820 177.875 102.990 ;
        RECT 176.850 101.600 177.310 102.650 ;
        RECT 177.480 101.460 177.650 102.820 ;
        RECT 178.045 102.560 178.510 102.950 ;
        RECT 177.820 101.750 178.170 102.370 ;
        RECT 178.340 101.970 178.510 102.560 ;
        RECT 178.680 102.340 178.850 103.120 ;
        RECT 179.020 103.020 179.190 103.360 ;
        RECT 179.425 103.190 179.755 103.620 ;
        RECT 179.925 103.020 180.095 103.360 ;
        RECT 180.390 103.160 180.760 103.620 ;
        RECT 179.020 102.850 180.095 103.020 ;
        RECT 180.930 102.990 181.100 103.450 ;
        RECT 181.335 103.110 182.205 103.450 ;
        RECT 182.375 103.160 182.625 103.620 ;
        RECT 180.540 102.820 181.100 102.990 ;
        RECT 180.540 102.680 180.710 102.820 ;
        RECT 179.210 102.510 180.710 102.680 ;
        RECT 181.405 102.650 181.865 102.940 ;
        RECT 178.680 102.170 180.370 102.340 ;
        RECT 178.340 101.750 178.695 101.970 ;
        RECT 178.865 101.460 179.035 102.170 ;
        RECT 179.240 101.750 180.030 102.000 ;
        RECT 180.200 101.990 180.370 102.170 ;
        RECT 180.540 101.820 180.710 102.510 ;
        RECT 176.980 101.070 177.310 101.430 ;
        RECT 177.480 101.290 177.975 101.460 ;
        RECT 178.180 101.290 179.035 101.460 ;
        RECT 179.910 101.070 180.240 101.530 ;
        RECT 180.450 101.430 180.710 101.820 ;
        RECT 180.900 102.640 181.865 102.650 ;
        RECT 182.035 102.730 182.205 103.110 ;
        RECT 182.795 103.070 182.965 103.360 ;
        RECT 183.145 103.240 183.475 103.620 ;
        RECT 182.795 102.900 183.595 103.070 ;
        RECT 180.900 102.480 181.575 102.640 ;
        RECT 182.035 102.560 183.255 102.730 ;
        RECT 180.900 101.690 181.110 102.480 ;
        RECT 182.035 102.470 182.205 102.560 ;
        RECT 181.280 101.690 181.630 102.310 ;
        RECT 181.800 102.300 182.205 102.470 ;
        RECT 181.800 101.520 181.970 102.300 ;
        RECT 182.140 101.850 182.360 102.130 ;
        RECT 182.540 102.020 183.080 102.390 ;
        RECT 183.425 102.310 183.595 102.900 ;
        RECT 183.815 102.480 184.120 103.620 ;
        RECT 184.290 102.430 184.545 103.310 ;
        RECT 185.730 102.690 185.900 103.450 ;
        RECT 186.115 102.860 186.445 103.620 ;
        RECT 185.730 102.520 186.445 102.690 ;
        RECT 186.615 102.545 186.870 103.450 ;
        RECT 183.425 102.280 184.165 102.310 ;
        RECT 182.140 101.680 182.670 101.850 ;
        RECT 180.450 101.260 180.800 101.430 ;
        RECT 181.020 101.240 181.970 101.520 ;
        RECT 182.140 101.070 182.330 101.510 ;
        RECT 182.500 101.450 182.670 101.680 ;
        RECT 182.840 101.620 183.080 102.020 ;
        RECT 183.250 101.980 184.165 102.280 ;
        RECT 183.250 101.805 183.575 101.980 ;
        RECT 183.250 101.450 183.570 101.805 ;
        RECT 184.335 101.780 184.545 102.430 ;
        RECT 185.640 101.970 185.995 102.340 ;
        RECT 186.275 102.310 186.445 102.520 ;
        RECT 186.275 101.980 186.530 102.310 ;
        RECT 186.275 101.790 186.445 101.980 ;
        RECT 186.700 101.815 186.870 102.545 ;
        RECT 187.045 102.470 187.305 103.620 ;
        RECT 187.485 102.950 187.740 103.450 ;
        RECT 187.910 103.120 188.240 103.620 ;
        RECT 187.485 102.780 188.235 102.950 ;
        RECT 187.485 101.960 187.835 102.610 ;
        RECT 182.500 101.280 183.570 101.450 ;
        RECT 183.815 101.070 184.120 101.530 ;
        RECT 184.290 101.250 184.545 101.780 ;
        RECT 185.730 101.620 186.445 101.790 ;
        RECT 185.730 101.240 185.900 101.620 ;
        RECT 186.115 101.070 186.445 101.450 ;
        RECT 186.615 101.240 186.870 101.815 ;
        RECT 187.045 101.070 187.305 101.910 ;
        RECT 188.005 101.790 188.235 102.780 ;
        RECT 187.485 101.620 188.235 101.790 ;
        RECT 187.485 101.330 187.740 101.620 ;
        RECT 187.910 101.070 188.240 101.450 ;
        RECT 188.410 101.330 188.580 103.450 ;
        RECT 188.750 102.650 189.075 103.435 ;
        RECT 189.245 103.160 189.495 103.620 ;
        RECT 189.665 103.120 189.915 103.450 ;
        RECT 190.130 103.120 190.810 103.450 ;
        RECT 189.665 102.990 189.835 103.120 ;
        RECT 189.440 102.820 189.835 102.990 ;
        RECT 188.810 101.600 189.270 102.650 ;
        RECT 189.440 101.460 189.610 102.820 ;
        RECT 190.005 102.560 190.470 102.950 ;
        RECT 189.780 101.750 190.130 102.370 ;
        RECT 190.300 101.970 190.470 102.560 ;
        RECT 190.640 102.340 190.810 103.120 ;
        RECT 190.980 103.020 191.150 103.360 ;
        RECT 191.385 103.190 191.715 103.620 ;
        RECT 191.885 103.020 192.055 103.360 ;
        RECT 192.350 103.160 192.720 103.620 ;
        RECT 190.980 102.850 192.055 103.020 ;
        RECT 192.890 102.990 193.060 103.450 ;
        RECT 193.295 103.110 194.165 103.450 ;
        RECT 194.335 103.160 194.585 103.620 ;
        RECT 192.500 102.820 193.060 102.990 ;
        RECT 192.500 102.680 192.670 102.820 ;
        RECT 191.170 102.510 192.670 102.680 ;
        RECT 193.365 102.650 193.825 102.940 ;
        RECT 190.640 102.170 192.330 102.340 ;
        RECT 190.300 101.750 190.655 101.970 ;
        RECT 190.825 101.460 190.995 102.170 ;
        RECT 191.200 101.750 191.990 102.000 ;
        RECT 192.160 101.990 192.330 102.170 ;
        RECT 192.500 101.820 192.670 102.510 ;
        RECT 188.940 101.070 189.270 101.430 ;
        RECT 189.440 101.290 189.935 101.460 ;
        RECT 190.140 101.290 190.995 101.460 ;
        RECT 191.870 101.070 192.200 101.530 ;
        RECT 192.410 101.430 192.670 101.820 ;
        RECT 192.860 102.640 193.825 102.650 ;
        RECT 193.995 102.730 194.165 103.110 ;
        RECT 194.755 103.070 194.925 103.360 ;
        RECT 195.105 103.240 195.435 103.620 ;
        RECT 194.755 102.900 195.555 103.070 ;
        RECT 192.860 102.480 193.535 102.640 ;
        RECT 193.995 102.560 195.215 102.730 ;
        RECT 192.860 101.690 193.070 102.480 ;
        RECT 193.995 102.470 194.165 102.560 ;
        RECT 193.240 101.690 193.590 102.310 ;
        RECT 193.760 102.300 194.165 102.470 ;
        RECT 193.760 101.520 193.930 102.300 ;
        RECT 194.100 101.850 194.320 102.130 ;
        RECT 194.500 102.020 195.040 102.390 ;
        RECT 195.385 102.310 195.555 102.900 ;
        RECT 195.775 102.480 196.080 103.620 ;
        RECT 196.250 102.430 196.505 103.310 ;
        RECT 196.685 102.470 196.945 103.620 ;
        RECT 197.120 102.545 197.375 103.450 ;
        RECT 197.545 102.860 197.875 103.620 ;
        RECT 198.090 102.690 198.260 103.450 ;
        RECT 195.385 102.280 196.125 102.310 ;
        RECT 194.100 101.680 194.630 101.850 ;
        RECT 192.410 101.260 192.760 101.430 ;
        RECT 192.980 101.240 193.930 101.520 ;
        RECT 194.100 101.070 194.290 101.510 ;
        RECT 194.460 101.450 194.630 101.680 ;
        RECT 194.800 101.620 195.040 102.020 ;
        RECT 195.210 101.980 196.125 102.280 ;
        RECT 195.210 101.805 195.535 101.980 ;
        RECT 195.210 101.450 195.530 101.805 ;
        RECT 196.295 101.780 196.505 102.430 ;
        RECT 194.460 101.280 195.530 101.450 ;
        RECT 195.775 101.070 196.080 101.530 ;
        RECT 196.250 101.250 196.505 101.780 ;
        RECT 196.685 101.070 196.945 101.910 ;
        RECT 197.120 101.815 197.290 102.545 ;
        RECT 197.545 102.520 198.260 102.690 ;
        RECT 197.545 102.310 197.715 102.520 ;
        RECT 198.985 102.470 199.245 103.620 ;
        RECT 199.420 102.545 199.675 103.450 ;
        RECT 199.845 102.860 200.175 103.620 ;
        RECT 200.390 102.690 200.560 103.450 ;
        RECT 197.460 101.980 197.715 102.310 ;
        RECT 197.120 101.240 197.375 101.815 ;
        RECT 197.545 101.790 197.715 101.980 ;
        RECT 197.995 101.970 198.350 102.340 ;
        RECT 197.545 101.620 198.260 101.790 ;
        RECT 197.545 101.070 197.875 101.450 ;
        RECT 198.090 101.240 198.260 101.620 ;
        RECT 198.985 101.070 199.245 101.910 ;
        RECT 199.420 101.815 199.590 102.545 ;
        RECT 199.845 102.520 200.560 102.690 ;
        RECT 199.845 102.310 200.015 102.520 ;
        RECT 200.820 102.455 201.110 103.620 ;
        RECT 201.285 102.470 201.545 103.620 ;
        RECT 201.720 102.545 201.975 103.450 ;
        RECT 202.145 102.860 202.475 103.620 ;
        RECT 202.690 102.690 202.860 103.450 ;
        RECT 203.585 102.950 203.840 103.450 ;
        RECT 204.010 103.120 204.340 103.620 ;
        RECT 203.585 102.780 204.335 102.950 ;
        RECT 199.760 101.980 200.015 102.310 ;
        RECT 199.420 101.240 199.675 101.815 ;
        RECT 199.845 101.790 200.015 101.980 ;
        RECT 200.295 101.970 200.650 102.340 ;
        RECT 199.845 101.620 200.560 101.790 ;
        RECT 199.845 101.070 200.175 101.450 ;
        RECT 200.390 101.240 200.560 101.620 ;
        RECT 200.820 101.070 201.110 101.795 ;
        RECT 201.285 101.070 201.545 101.910 ;
        RECT 201.720 101.815 201.890 102.545 ;
        RECT 202.145 102.520 202.860 102.690 ;
        RECT 202.145 102.310 202.315 102.520 ;
        RECT 202.060 101.980 202.315 102.310 ;
        RECT 201.720 101.240 201.975 101.815 ;
        RECT 202.145 101.790 202.315 101.980 ;
        RECT 202.595 101.970 202.950 102.340 ;
        RECT 203.585 101.960 203.935 102.610 ;
        RECT 204.105 101.790 204.335 102.780 ;
        RECT 202.145 101.620 202.860 101.790 ;
        RECT 202.145 101.070 202.475 101.450 ;
        RECT 202.690 101.240 202.860 101.620 ;
        RECT 203.585 101.620 204.335 101.790 ;
        RECT 203.585 101.330 203.840 101.620 ;
        RECT 204.010 101.070 204.340 101.450 ;
        RECT 204.510 101.330 204.680 103.450 ;
        RECT 204.850 102.650 205.175 103.435 ;
        RECT 205.345 103.160 205.595 103.620 ;
        RECT 205.765 103.120 206.015 103.450 ;
        RECT 206.230 103.120 206.910 103.450 ;
        RECT 205.765 102.990 205.935 103.120 ;
        RECT 205.540 102.820 205.935 102.990 ;
        RECT 204.910 101.600 205.370 102.650 ;
        RECT 205.540 101.460 205.710 102.820 ;
        RECT 206.105 102.560 206.570 102.950 ;
        RECT 205.880 101.750 206.230 102.370 ;
        RECT 206.400 101.970 206.570 102.560 ;
        RECT 206.740 102.340 206.910 103.120 ;
        RECT 207.080 103.020 207.250 103.360 ;
        RECT 207.485 103.190 207.815 103.620 ;
        RECT 207.985 103.020 208.155 103.360 ;
        RECT 208.450 103.160 208.820 103.620 ;
        RECT 207.080 102.850 208.155 103.020 ;
        RECT 208.990 102.990 209.160 103.450 ;
        RECT 209.395 103.110 210.265 103.450 ;
        RECT 210.435 103.160 210.685 103.620 ;
        RECT 208.600 102.820 209.160 102.990 ;
        RECT 208.600 102.680 208.770 102.820 ;
        RECT 207.270 102.510 208.770 102.680 ;
        RECT 209.465 102.650 209.925 102.940 ;
        RECT 206.740 102.170 208.430 102.340 ;
        RECT 206.400 101.750 206.755 101.970 ;
        RECT 206.925 101.460 207.095 102.170 ;
        RECT 207.300 101.750 208.090 102.000 ;
        RECT 208.260 101.990 208.430 102.170 ;
        RECT 208.600 101.820 208.770 102.510 ;
        RECT 205.040 101.070 205.370 101.430 ;
        RECT 205.540 101.290 206.035 101.460 ;
        RECT 206.240 101.290 207.095 101.460 ;
        RECT 207.970 101.070 208.300 101.530 ;
        RECT 208.510 101.430 208.770 101.820 ;
        RECT 208.960 102.640 209.925 102.650 ;
        RECT 210.095 102.730 210.265 103.110 ;
        RECT 210.855 103.070 211.025 103.360 ;
        RECT 211.205 103.240 211.535 103.620 ;
        RECT 210.855 102.900 211.655 103.070 ;
        RECT 208.960 102.480 209.635 102.640 ;
        RECT 210.095 102.560 211.315 102.730 ;
        RECT 208.960 101.690 209.170 102.480 ;
        RECT 210.095 102.470 210.265 102.560 ;
        RECT 209.340 101.690 209.690 102.310 ;
        RECT 209.860 102.300 210.265 102.470 ;
        RECT 209.860 101.520 210.030 102.300 ;
        RECT 210.200 101.850 210.420 102.130 ;
        RECT 210.600 102.020 211.140 102.390 ;
        RECT 211.485 102.310 211.655 102.900 ;
        RECT 211.875 102.480 212.180 103.620 ;
        RECT 212.350 102.430 212.605 103.310 ;
        RECT 211.485 102.280 212.225 102.310 ;
        RECT 210.200 101.680 210.730 101.850 ;
        RECT 208.510 101.260 208.860 101.430 ;
        RECT 209.080 101.240 210.030 101.520 ;
        RECT 210.200 101.070 210.390 101.510 ;
        RECT 210.560 101.450 210.730 101.680 ;
        RECT 210.900 101.620 211.140 102.020 ;
        RECT 211.310 101.980 212.225 102.280 ;
        RECT 211.310 101.805 211.635 101.980 ;
        RECT 211.310 101.450 211.630 101.805 ;
        RECT 212.395 101.780 212.605 102.430 ;
        RECT 210.560 101.280 211.630 101.450 ;
        RECT 211.875 101.070 212.180 101.530 ;
        RECT 212.350 101.250 212.605 101.780 ;
        RECT 212.785 102.480 213.120 103.450 ;
        RECT 213.290 102.480 213.460 103.620 ;
        RECT 213.630 103.280 215.660 103.450 ;
        RECT 212.785 101.810 212.955 102.480 ;
        RECT 213.630 102.310 213.800 103.280 ;
        RECT 213.125 101.980 213.380 102.310 ;
        RECT 213.605 101.980 213.800 102.310 ;
        RECT 213.970 102.940 215.095 103.110 ;
        RECT 213.210 101.810 213.380 101.980 ;
        RECT 213.970 101.810 214.140 102.940 ;
        RECT 212.785 101.240 213.040 101.810 ;
        RECT 213.210 101.640 214.140 101.810 ;
        RECT 214.310 102.600 215.320 102.770 ;
        RECT 214.310 101.800 214.480 102.600 ;
        RECT 213.965 101.605 214.140 101.640 ;
        RECT 213.210 101.070 213.540 101.470 ;
        RECT 213.965 101.240 214.495 101.605 ;
        RECT 214.685 101.580 214.960 102.400 ;
        RECT 214.680 101.410 214.960 101.580 ;
        RECT 214.685 101.240 214.960 101.410 ;
        RECT 215.130 101.240 215.320 102.600 ;
        RECT 215.490 102.615 215.660 103.280 ;
        RECT 215.830 102.860 216.000 103.620 ;
        RECT 216.235 102.860 216.750 103.270 ;
        RECT 215.490 102.425 216.240 102.615 ;
        RECT 216.410 102.050 216.750 102.860 ;
        RECT 215.520 101.880 216.750 102.050 ;
        RECT 217.385 102.430 217.640 103.310 ;
        RECT 217.810 102.480 218.115 103.620 ;
        RECT 218.455 103.240 218.785 103.620 ;
        RECT 218.965 103.070 219.135 103.360 ;
        RECT 219.305 103.160 219.555 103.620 ;
        RECT 218.335 102.900 219.135 103.070 ;
        RECT 219.725 103.110 220.595 103.450 ;
        RECT 215.500 101.070 216.010 101.605 ;
        RECT 216.230 101.275 216.475 101.880 ;
        RECT 217.385 101.780 217.595 102.430 ;
        RECT 218.335 102.310 218.505 102.900 ;
        RECT 219.725 102.730 219.895 103.110 ;
        RECT 220.830 102.990 221.000 103.450 ;
        RECT 221.170 103.160 221.540 103.620 ;
        RECT 221.835 103.020 222.005 103.360 ;
        RECT 222.175 103.190 222.505 103.620 ;
        RECT 222.740 103.020 222.910 103.360 ;
        RECT 218.675 102.560 219.895 102.730 ;
        RECT 220.065 102.650 220.525 102.940 ;
        RECT 220.830 102.820 221.390 102.990 ;
        RECT 221.835 102.850 222.910 103.020 ;
        RECT 223.080 103.120 223.760 103.450 ;
        RECT 223.975 103.120 224.225 103.450 ;
        RECT 224.395 103.160 224.645 103.620 ;
        RECT 221.220 102.680 221.390 102.820 ;
        RECT 220.065 102.640 221.030 102.650 ;
        RECT 219.725 102.470 219.895 102.560 ;
        RECT 220.355 102.480 221.030 102.640 ;
        RECT 217.765 102.280 218.505 102.310 ;
        RECT 217.765 101.980 218.680 102.280 ;
        RECT 218.355 101.805 218.680 101.980 ;
        RECT 217.385 101.250 217.640 101.780 ;
        RECT 217.810 101.070 218.115 101.530 ;
        RECT 218.360 101.450 218.680 101.805 ;
        RECT 218.850 102.020 219.390 102.390 ;
        RECT 219.725 102.300 220.130 102.470 ;
        RECT 218.850 101.620 219.090 102.020 ;
        RECT 219.570 101.850 219.790 102.130 ;
        RECT 219.260 101.680 219.790 101.850 ;
        RECT 219.260 101.450 219.430 101.680 ;
        RECT 219.960 101.520 220.130 102.300 ;
        RECT 220.300 101.690 220.650 102.310 ;
        RECT 220.820 101.690 221.030 102.480 ;
        RECT 221.220 102.510 222.720 102.680 ;
        RECT 221.220 101.820 221.390 102.510 ;
        RECT 223.080 102.340 223.250 103.120 ;
        RECT 224.055 102.990 224.225 103.120 ;
        RECT 221.560 102.170 223.250 102.340 ;
        RECT 223.420 102.560 223.885 102.950 ;
        RECT 224.055 102.820 224.450 102.990 ;
        RECT 221.560 101.990 221.730 102.170 ;
        RECT 218.360 101.280 219.430 101.450 ;
        RECT 219.600 101.070 219.790 101.510 ;
        RECT 219.960 101.240 220.910 101.520 ;
        RECT 221.220 101.430 221.480 101.820 ;
        RECT 221.900 101.750 222.690 102.000 ;
        RECT 221.130 101.260 221.480 101.430 ;
        RECT 221.690 101.070 222.020 101.530 ;
        RECT 222.895 101.460 223.065 102.170 ;
        RECT 223.420 101.970 223.590 102.560 ;
        RECT 223.235 101.750 223.590 101.970 ;
        RECT 223.760 101.750 224.110 102.370 ;
        RECT 224.280 101.460 224.450 102.820 ;
        RECT 224.815 102.650 225.140 103.435 ;
        RECT 224.620 101.600 225.080 102.650 ;
        RECT 222.895 101.290 223.750 101.460 ;
        RECT 223.955 101.290 224.450 101.460 ;
        RECT 224.620 101.070 224.950 101.430 ;
        RECT 225.310 101.330 225.480 103.450 ;
        RECT 225.650 103.120 225.980 103.620 ;
        RECT 226.150 102.950 226.405 103.450 ;
        RECT 225.655 102.780 226.405 102.950 ;
        RECT 225.655 101.790 225.885 102.780 ;
        RECT 226.055 101.960 226.405 102.610 ;
        RECT 226.580 102.455 226.870 103.620 ;
        RECT 227.045 102.480 227.380 103.450 ;
        RECT 227.550 102.480 227.720 103.620 ;
        RECT 227.890 103.280 229.920 103.450 ;
        RECT 227.045 101.810 227.215 102.480 ;
        RECT 227.890 102.310 228.060 103.280 ;
        RECT 227.385 101.980 227.640 102.310 ;
        RECT 227.865 101.980 228.060 102.310 ;
        RECT 228.230 102.940 229.355 103.110 ;
        RECT 227.470 101.810 227.640 101.980 ;
        RECT 228.230 101.810 228.400 102.940 ;
        RECT 225.655 101.620 226.405 101.790 ;
        RECT 225.650 101.070 225.980 101.450 ;
        RECT 226.150 101.330 226.405 101.620 ;
        RECT 226.580 101.070 226.870 101.795 ;
        RECT 227.045 101.240 227.300 101.810 ;
        RECT 227.470 101.640 228.400 101.810 ;
        RECT 228.570 102.600 229.580 102.770 ;
        RECT 228.570 101.800 228.740 102.600 ;
        RECT 228.225 101.605 228.400 101.640 ;
        RECT 227.470 101.070 227.800 101.470 ;
        RECT 228.225 101.240 228.755 101.605 ;
        RECT 228.945 101.580 229.220 102.400 ;
        RECT 228.940 101.410 229.220 101.580 ;
        RECT 228.945 101.240 229.220 101.410 ;
        RECT 229.390 101.240 229.580 102.600 ;
        RECT 229.750 102.615 229.920 103.280 ;
        RECT 230.090 102.860 230.260 103.620 ;
        RECT 230.495 102.860 231.010 103.270 ;
        RECT 229.750 102.425 230.500 102.615 ;
        RECT 230.670 102.050 231.010 102.860 ;
        RECT 231.185 102.470 231.445 103.620 ;
        RECT 231.620 102.545 231.875 103.450 ;
        RECT 232.045 102.860 232.375 103.620 ;
        RECT 232.590 102.690 232.760 103.450 ;
        RECT 229.780 101.880 231.010 102.050 ;
        RECT 229.760 101.070 230.270 101.605 ;
        RECT 230.490 101.275 230.735 101.880 ;
        RECT 231.185 101.070 231.445 101.910 ;
        RECT 231.620 101.815 231.790 102.545 ;
        RECT 232.045 102.520 232.760 102.690 ;
        RECT 233.020 102.530 236.530 103.620 ;
        RECT 237.165 102.950 237.420 103.450 ;
        RECT 237.590 103.120 237.920 103.620 ;
        RECT 237.165 102.780 237.915 102.950 ;
        RECT 232.045 102.310 232.215 102.520 ;
        RECT 231.960 101.980 232.215 102.310 ;
        RECT 231.620 101.240 231.875 101.815 ;
        RECT 232.045 101.790 232.215 101.980 ;
        RECT 232.495 101.970 232.850 102.340 ;
        RECT 233.020 101.840 234.670 102.360 ;
        RECT 234.840 102.010 236.530 102.530 ;
        RECT 237.165 101.960 237.515 102.610 ;
        RECT 232.045 101.620 232.760 101.790 ;
        RECT 232.045 101.070 232.375 101.450 ;
        RECT 232.590 101.240 232.760 101.620 ;
        RECT 233.020 101.070 236.530 101.840 ;
        RECT 237.685 101.790 237.915 102.780 ;
        RECT 237.165 101.620 237.915 101.790 ;
        RECT 237.165 101.330 237.420 101.620 ;
        RECT 237.590 101.070 237.920 101.450 ;
        RECT 238.090 101.330 238.260 103.450 ;
        RECT 238.430 102.650 238.755 103.435 ;
        RECT 238.925 103.160 239.175 103.620 ;
        RECT 239.345 103.120 239.595 103.450 ;
        RECT 239.810 103.120 240.490 103.450 ;
        RECT 239.345 102.990 239.515 103.120 ;
        RECT 239.120 102.820 239.515 102.990 ;
        RECT 238.490 101.600 238.950 102.650 ;
        RECT 239.120 101.460 239.290 102.820 ;
        RECT 239.685 102.560 240.150 102.950 ;
        RECT 239.460 101.750 239.810 102.370 ;
        RECT 239.980 101.970 240.150 102.560 ;
        RECT 240.320 102.340 240.490 103.120 ;
        RECT 240.660 103.020 240.830 103.360 ;
        RECT 241.065 103.190 241.395 103.620 ;
        RECT 241.565 103.020 241.735 103.360 ;
        RECT 242.030 103.160 242.400 103.620 ;
        RECT 240.660 102.850 241.735 103.020 ;
        RECT 242.570 102.990 242.740 103.450 ;
        RECT 242.975 103.110 243.845 103.450 ;
        RECT 244.015 103.160 244.265 103.620 ;
        RECT 242.180 102.820 242.740 102.990 ;
        RECT 242.180 102.680 242.350 102.820 ;
        RECT 240.850 102.510 242.350 102.680 ;
        RECT 243.045 102.650 243.505 102.940 ;
        RECT 240.320 102.170 242.010 102.340 ;
        RECT 239.980 101.750 240.335 101.970 ;
        RECT 240.505 101.460 240.675 102.170 ;
        RECT 240.880 101.750 241.670 102.000 ;
        RECT 241.840 101.990 242.010 102.170 ;
        RECT 242.180 101.820 242.350 102.510 ;
        RECT 238.620 101.070 238.950 101.430 ;
        RECT 239.120 101.290 239.615 101.460 ;
        RECT 239.820 101.290 240.675 101.460 ;
        RECT 241.550 101.070 241.880 101.530 ;
        RECT 242.090 101.430 242.350 101.820 ;
        RECT 242.540 102.640 243.505 102.650 ;
        RECT 243.675 102.730 243.845 103.110 ;
        RECT 244.435 103.070 244.605 103.360 ;
        RECT 244.785 103.240 245.115 103.620 ;
        RECT 244.435 102.900 245.235 103.070 ;
        RECT 242.540 102.480 243.215 102.640 ;
        RECT 243.675 102.560 244.895 102.730 ;
        RECT 242.540 101.690 242.750 102.480 ;
        RECT 243.675 102.470 243.845 102.560 ;
        RECT 242.920 101.690 243.270 102.310 ;
        RECT 243.440 102.300 243.845 102.470 ;
        RECT 243.440 101.520 243.610 102.300 ;
        RECT 243.780 101.850 244.000 102.130 ;
        RECT 244.180 102.020 244.720 102.390 ;
        RECT 245.065 102.310 245.235 102.900 ;
        RECT 245.455 102.480 245.760 103.620 ;
        RECT 245.930 102.430 246.185 103.310 ;
        RECT 245.065 102.280 245.805 102.310 ;
        RECT 243.780 101.680 244.310 101.850 ;
        RECT 242.090 101.260 242.440 101.430 ;
        RECT 242.660 101.240 243.610 101.520 ;
        RECT 243.780 101.070 243.970 101.510 ;
        RECT 244.140 101.450 244.310 101.680 ;
        RECT 244.480 101.620 244.720 102.020 ;
        RECT 244.890 101.980 245.805 102.280 ;
        RECT 244.890 101.805 245.215 101.980 ;
        RECT 244.890 101.450 245.210 101.805 ;
        RECT 245.975 101.780 246.185 102.430 ;
        RECT 244.140 101.280 245.210 101.450 ;
        RECT 245.455 101.070 245.760 101.530 ;
        RECT 245.930 101.250 246.185 101.780 ;
        RECT 246.365 102.480 246.700 103.450 ;
        RECT 246.870 102.480 247.040 103.620 ;
        RECT 247.210 103.280 249.240 103.450 ;
        RECT 246.365 101.810 246.535 102.480 ;
        RECT 247.210 102.310 247.380 103.280 ;
        RECT 246.705 101.980 246.960 102.310 ;
        RECT 247.185 101.980 247.380 102.310 ;
        RECT 247.550 102.940 248.675 103.110 ;
        RECT 246.790 101.810 246.960 101.980 ;
        RECT 247.550 101.810 247.720 102.940 ;
        RECT 246.365 101.240 246.620 101.810 ;
        RECT 246.790 101.640 247.720 101.810 ;
        RECT 247.890 102.600 248.900 102.770 ;
        RECT 247.890 101.800 248.060 102.600 ;
        RECT 247.545 101.605 247.720 101.640 ;
        RECT 246.790 101.070 247.120 101.470 ;
        RECT 247.545 101.240 248.075 101.605 ;
        RECT 248.265 101.580 248.540 102.400 ;
        RECT 248.260 101.410 248.540 101.580 ;
        RECT 248.265 101.240 248.540 101.410 ;
        RECT 248.710 101.240 248.900 102.600 ;
        RECT 249.070 102.615 249.240 103.280 ;
        RECT 249.410 102.860 249.580 103.620 ;
        RECT 249.815 102.860 250.330 103.270 ;
        RECT 249.070 102.425 249.820 102.615 ;
        RECT 249.990 102.050 250.330 102.860 ;
        RECT 250.590 102.690 250.760 103.450 ;
        RECT 250.975 102.860 251.305 103.620 ;
        RECT 250.590 102.520 251.305 102.690 ;
        RECT 251.475 102.545 251.730 103.450 ;
        RECT 249.100 101.880 250.330 102.050 ;
        RECT 250.500 101.970 250.855 102.340 ;
        RECT 251.135 102.310 251.305 102.520 ;
        RECT 251.135 101.980 251.390 102.310 ;
        RECT 249.080 101.070 249.590 101.605 ;
        RECT 249.810 101.275 250.055 101.880 ;
        RECT 251.135 101.790 251.305 101.980 ;
        RECT 251.560 101.815 251.730 102.545 ;
        RECT 251.905 102.470 252.165 103.620 ;
        RECT 252.340 102.455 252.630 103.620 ;
        RECT 252.805 102.480 253.140 103.450 ;
        RECT 253.310 102.480 253.480 103.620 ;
        RECT 253.650 103.280 255.680 103.450 ;
        RECT 250.590 101.620 251.305 101.790 ;
        RECT 250.590 101.240 250.760 101.620 ;
        RECT 250.975 101.070 251.305 101.450 ;
        RECT 251.475 101.240 251.730 101.815 ;
        RECT 251.905 101.070 252.165 101.910 ;
        RECT 252.805 101.810 252.975 102.480 ;
        RECT 253.650 102.310 253.820 103.280 ;
        RECT 253.145 101.980 253.400 102.310 ;
        RECT 253.625 101.980 253.820 102.310 ;
        RECT 253.990 102.940 255.115 103.110 ;
        RECT 253.230 101.810 253.400 101.980 ;
        RECT 253.990 101.810 254.160 102.940 ;
        RECT 252.340 101.070 252.630 101.795 ;
        RECT 252.805 101.240 253.060 101.810 ;
        RECT 253.230 101.640 254.160 101.810 ;
        RECT 254.330 102.600 255.340 102.770 ;
        RECT 254.330 101.800 254.500 102.600 ;
        RECT 254.705 102.260 254.980 102.400 ;
        RECT 254.700 102.090 254.980 102.260 ;
        RECT 253.985 101.605 254.160 101.640 ;
        RECT 253.230 101.070 253.560 101.470 ;
        RECT 253.985 101.240 254.515 101.605 ;
        RECT 254.705 101.240 254.980 102.090 ;
        RECT 255.150 101.240 255.340 102.600 ;
        RECT 255.510 102.615 255.680 103.280 ;
        RECT 255.850 102.860 256.020 103.620 ;
        RECT 256.255 102.860 256.770 103.270 ;
        RECT 255.510 102.425 256.260 102.615 ;
        RECT 256.430 102.050 256.770 102.860 ;
        RECT 257.405 102.950 257.660 103.450 ;
        RECT 257.830 103.120 258.160 103.620 ;
        RECT 257.405 102.780 258.155 102.950 ;
        RECT 255.540 101.880 256.770 102.050 ;
        RECT 257.405 101.960 257.755 102.610 ;
        RECT 255.520 101.070 256.030 101.605 ;
        RECT 256.250 101.275 256.495 101.880 ;
        RECT 257.925 101.790 258.155 102.780 ;
        RECT 257.405 101.620 258.155 101.790 ;
        RECT 257.405 101.330 257.660 101.620 ;
        RECT 257.830 101.070 258.160 101.450 ;
        RECT 258.330 101.330 258.500 103.450 ;
        RECT 258.670 102.650 258.995 103.435 ;
        RECT 259.165 103.160 259.415 103.620 ;
        RECT 259.585 103.120 259.835 103.450 ;
        RECT 260.050 103.120 260.730 103.450 ;
        RECT 259.585 102.990 259.755 103.120 ;
        RECT 259.360 102.820 259.755 102.990 ;
        RECT 258.730 101.600 259.190 102.650 ;
        RECT 259.360 101.460 259.530 102.820 ;
        RECT 259.925 102.560 260.390 102.950 ;
        RECT 259.700 101.750 260.050 102.370 ;
        RECT 260.220 101.970 260.390 102.560 ;
        RECT 260.560 102.340 260.730 103.120 ;
        RECT 260.900 103.020 261.070 103.360 ;
        RECT 261.305 103.190 261.635 103.620 ;
        RECT 261.805 103.020 261.975 103.360 ;
        RECT 262.270 103.160 262.640 103.620 ;
        RECT 260.900 102.850 261.975 103.020 ;
        RECT 262.810 102.990 262.980 103.450 ;
        RECT 263.215 103.110 264.085 103.450 ;
        RECT 264.255 103.160 264.505 103.620 ;
        RECT 262.420 102.820 262.980 102.990 ;
        RECT 262.420 102.680 262.590 102.820 ;
        RECT 261.090 102.510 262.590 102.680 ;
        RECT 263.285 102.650 263.745 102.940 ;
        RECT 260.560 102.170 262.250 102.340 ;
        RECT 260.220 101.750 260.575 101.970 ;
        RECT 260.745 101.460 260.915 102.170 ;
        RECT 261.120 101.750 261.910 102.000 ;
        RECT 262.080 101.990 262.250 102.170 ;
        RECT 262.420 101.820 262.590 102.510 ;
        RECT 258.860 101.070 259.190 101.430 ;
        RECT 259.360 101.290 259.855 101.460 ;
        RECT 260.060 101.290 260.915 101.460 ;
        RECT 261.790 101.070 262.120 101.530 ;
        RECT 262.330 101.430 262.590 101.820 ;
        RECT 262.780 102.640 263.745 102.650 ;
        RECT 263.915 102.730 264.085 103.110 ;
        RECT 264.675 103.070 264.845 103.360 ;
        RECT 265.025 103.240 265.355 103.620 ;
        RECT 264.675 102.900 265.475 103.070 ;
        RECT 262.780 102.480 263.455 102.640 ;
        RECT 263.915 102.560 265.135 102.730 ;
        RECT 262.780 101.690 262.990 102.480 ;
        RECT 263.915 102.470 264.085 102.560 ;
        RECT 263.160 101.690 263.510 102.310 ;
        RECT 263.680 102.300 264.085 102.470 ;
        RECT 263.680 101.520 263.850 102.300 ;
        RECT 264.020 101.850 264.240 102.130 ;
        RECT 264.420 102.020 264.960 102.390 ;
        RECT 265.305 102.310 265.475 102.900 ;
        RECT 265.695 102.480 266.000 103.620 ;
        RECT 266.170 102.430 266.425 103.310 ;
        RECT 266.605 102.950 266.860 103.450 ;
        RECT 267.030 103.120 267.360 103.620 ;
        RECT 266.605 102.780 267.355 102.950 ;
        RECT 265.305 102.280 266.045 102.310 ;
        RECT 264.020 101.680 264.550 101.850 ;
        RECT 262.330 101.260 262.680 101.430 ;
        RECT 262.900 101.240 263.850 101.520 ;
        RECT 264.020 101.070 264.210 101.510 ;
        RECT 264.380 101.450 264.550 101.680 ;
        RECT 264.720 101.620 264.960 102.020 ;
        RECT 265.130 101.980 266.045 102.280 ;
        RECT 265.130 101.805 265.455 101.980 ;
        RECT 265.130 101.450 265.450 101.805 ;
        RECT 266.215 101.780 266.425 102.430 ;
        RECT 266.605 101.960 266.955 102.610 ;
        RECT 267.125 101.790 267.355 102.780 ;
        RECT 264.380 101.280 265.450 101.450 ;
        RECT 265.695 101.070 266.000 101.530 ;
        RECT 266.170 101.250 266.425 101.780 ;
        RECT 266.605 101.620 267.355 101.790 ;
        RECT 266.605 101.330 266.860 101.620 ;
        RECT 267.030 101.070 267.360 101.450 ;
        RECT 267.530 101.330 267.700 103.450 ;
        RECT 267.870 102.650 268.195 103.435 ;
        RECT 268.365 103.160 268.615 103.620 ;
        RECT 268.785 103.120 269.035 103.450 ;
        RECT 269.250 103.120 269.930 103.450 ;
        RECT 268.785 102.990 268.955 103.120 ;
        RECT 268.560 102.820 268.955 102.990 ;
        RECT 267.930 101.600 268.390 102.650 ;
        RECT 268.560 101.460 268.730 102.820 ;
        RECT 269.125 102.560 269.590 102.950 ;
        RECT 268.900 101.750 269.250 102.370 ;
        RECT 269.420 101.970 269.590 102.560 ;
        RECT 269.760 102.340 269.930 103.120 ;
        RECT 270.100 103.020 270.270 103.360 ;
        RECT 270.505 103.190 270.835 103.620 ;
        RECT 271.005 103.020 271.175 103.360 ;
        RECT 271.470 103.160 271.840 103.620 ;
        RECT 270.100 102.850 271.175 103.020 ;
        RECT 272.010 102.990 272.180 103.450 ;
        RECT 272.415 103.110 273.285 103.450 ;
        RECT 273.455 103.160 273.705 103.620 ;
        RECT 271.620 102.820 272.180 102.990 ;
        RECT 271.620 102.680 271.790 102.820 ;
        RECT 270.290 102.510 271.790 102.680 ;
        RECT 272.485 102.650 272.945 102.940 ;
        RECT 269.760 102.170 271.450 102.340 ;
        RECT 269.420 101.750 269.775 101.970 ;
        RECT 269.945 101.460 270.115 102.170 ;
        RECT 270.320 101.750 271.110 102.000 ;
        RECT 271.280 101.990 271.450 102.170 ;
        RECT 271.620 101.820 271.790 102.510 ;
        RECT 268.060 101.070 268.390 101.430 ;
        RECT 268.560 101.290 269.055 101.460 ;
        RECT 269.260 101.290 270.115 101.460 ;
        RECT 270.990 101.070 271.320 101.530 ;
        RECT 271.530 101.430 271.790 101.820 ;
        RECT 271.980 102.640 272.945 102.650 ;
        RECT 273.115 102.730 273.285 103.110 ;
        RECT 273.875 103.070 274.045 103.360 ;
        RECT 274.225 103.240 274.555 103.620 ;
        RECT 273.875 102.900 274.675 103.070 ;
        RECT 271.980 102.480 272.655 102.640 ;
        RECT 273.115 102.560 274.335 102.730 ;
        RECT 271.980 101.690 272.190 102.480 ;
        RECT 273.115 102.470 273.285 102.560 ;
        RECT 272.360 101.690 272.710 102.310 ;
        RECT 272.880 102.300 273.285 102.470 ;
        RECT 272.880 101.520 273.050 102.300 ;
        RECT 273.220 101.850 273.440 102.130 ;
        RECT 273.620 102.020 274.160 102.390 ;
        RECT 274.505 102.310 274.675 102.900 ;
        RECT 274.895 102.480 275.200 103.620 ;
        RECT 275.370 102.430 275.625 103.310 ;
        RECT 275.805 102.470 276.065 103.620 ;
        RECT 276.240 102.545 276.495 103.450 ;
        RECT 276.665 102.860 276.995 103.620 ;
        RECT 277.210 102.690 277.380 103.450 ;
        RECT 274.505 102.280 275.245 102.310 ;
        RECT 273.220 101.680 273.750 101.850 ;
        RECT 271.530 101.260 271.880 101.430 ;
        RECT 272.100 101.240 273.050 101.520 ;
        RECT 273.220 101.070 273.410 101.510 ;
        RECT 273.580 101.450 273.750 101.680 ;
        RECT 273.920 101.620 274.160 102.020 ;
        RECT 274.330 101.980 275.245 102.280 ;
        RECT 274.330 101.805 274.655 101.980 ;
        RECT 274.330 101.450 274.650 101.805 ;
        RECT 275.415 101.780 275.625 102.430 ;
        RECT 273.580 101.280 274.650 101.450 ;
        RECT 274.895 101.070 275.200 101.530 ;
        RECT 275.370 101.250 275.625 101.780 ;
        RECT 275.805 101.070 276.065 101.910 ;
        RECT 276.240 101.815 276.410 102.545 ;
        RECT 276.665 102.520 277.380 102.690 ;
        RECT 276.665 102.310 276.835 102.520 ;
        RECT 278.100 102.455 278.390 103.620 ;
        RECT 278.565 102.430 278.820 103.310 ;
        RECT 278.990 102.480 279.295 103.620 ;
        RECT 279.635 103.240 279.965 103.620 ;
        RECT 280.145 103.070 280.315 103.360 ;
        RECT 280.485 103.160 280.735 103.620 ;
        RECT 279.515 102.900 280.315 103.070 ;
        RECT 280.905 103.110 281.775 103.450 ;
        RECT 276.580 101.980 276.835 102.310 ;
        RECT 276.240 101.240 276.495 101.815 ;
        RECT 276.665 101.790 276.835 101.980 ;
        RECT 277.115 101.970 277.470 102.340 ;
        RECT 276.665 101.620 277.380 101.790 ;
        RECT 276.665 101.070 276.995 101.450 ;
        RECT 277.210 101.240 277.380 101.620 ;
        RECT 278.100 101.070 278.390 101.795 ;
        RECT 278.565 101.780 278.775 102.430 ;
        RECT 279.515 102.310 279.685 102.900 ;
        RECT 280.905 102.730 281.075 103.110 ;
        RECT 282.010 102.990 282.180 103.450 ;
        RECT 282.350 103.160 282.720 103.620 ;
        RECT 283.015 103.020 283.185 103.360 ;
        RECT 283.355 103.190 283.685 103.620 ;
        RECT 283.920 103.020 284.090 103.360 ;
        RECT 279.855 102.560 281.075 102.730 ;
        RECT 281.245 102.650 281.705 102.940 ;
        RECT 282.010 102.820 282.570 102.990 ;
        RECT 283.015 102.850 284.090 103.020 ;
        RECT 284.260 103.120 284.940 103.450 ;
        RECT 285.155 103.120 285.405 103.450 ;
        RECT 285.575 103.160 285.825 103.620 ;
        RECT 282.400 102.680 282.570 102.820 ;
        RECT 281.245 102.640 282.210 102.650 ;
        RECT 280.905 102.470 281.075 102.560 ;
        RECT 281.535 102.480 282.210 102.640 ;
        RECT 278.945 102.280 279.685 102.310 ;
        RECT 278.945 101.980 279.860 102.280 ;
        RECT 279.535 101.805 279.860 101.980 ;
        RECT 278.565 101.250 278.820 101.780 ;
        RECT 278.990 101.070 279.295 101.530 ;
        RECT 279.540 101.450 279.860 101.805 ;
        RECT 280.030 102.020 280.570 102.390 ;
        RECT 280.905 102.300 281.310 102.470 ;
        RECT 280.030 101.620 280.270 102.020 ;
        RECT 280.750 101.850 280.970 102.130 ;
        RECT 280.440 101.680 280.970 101.850 ;
        RECT 280.440 101.450 280.610 101.680 ;
        RECT 281.140 101.520 281.310 102.300 ;
        RECT 281.480 101.690 281.830 102.310 ;
        RECT 282.000 101.690 282.210 102.480 ;
        RECT 282.400 102.510 283.900 102.680 ;
        RECT 282.400 101.820 282.570 102.510 ;
        RECT 284.260 102.340 284.430 103.120 ;
        RECT 285.235 102.990 285.405 103.120 ;
        RECT 282.740 102.170 284.430 102.340 ;
        RECT 284.600 102.560 285.065 102.950 ;
        RECT 285.235 102.820 285.630 102.990 ;
        RECT 282.740 101.990 282.910 102.170 ;
        RECT 279.540 101.280 280.610 101.450 ;
        RECT 280.780 101.070 280.970 101.510 ;
        RECT 281.140 101.240 282.090 101.520 ;
        RECT 282.400 101.430 282.660 101.820 ;
        RECT 283.080 101.750 283.870 102.000 ;
        RECT 282.310 101.260 282.660 101.430 ;
        RECT 282.870 101.070 283.200 101.530 ;
        RECT 284.075 101.460 284.245 102.170 ;
        RECT 284.600 101.970 284.770 102.560 ;
        RECT 284.415 101.750 284.770 101.970 ;
        RECT 284.940 101.750 285.290 102.370 ;
        RECT 285.460 101.460 285.630 102.820 ;
        RECT 285.995 102.650 286.320 103.435 ;
        RECT 285.800 101.600 286.260 102.650 ;
        RECT 284.075 101.290 284.930 101.460 ;
        RECT 285.135 101.290 285.630 101.460 ;
        RECT 285.800 101.070 286.130 101.430 ;
        RECT 286.490 101.330 286.660 103.450 ;
        RECT 286.830 103.120 287.160 103.620 ;
        RECT 287.330 102.950 287.585 103.450 ;
        RECT 286.835 102.780 287.585 102.950 ;
        RECT 286.835 101.790 287.065 102.780 ;
        RECT 287.235 101.960 287.585 102.610 ;
        RECT 287.765 102.430 288.020 103.310 ;
        RECT 288.190 102.480 288.495 103.620 ;
        RECT 288.835 103.240 289.165 103.620 ;
        RECT 289.345 103.070 289.515 103.360 ;
        RECT 289.685 103.160 289.935 103.620 ;
        RECT 288.715 102.900 289.515 103.070 ;
        RECT 290.105 103.110 290.975 103.450 ;
        RECT 286.835 101.620 287.585 101.790 ;
        RECT 286.830 101.070 287.160 101.450 ;
        RECT 287.330 101.330 287.585 101.620 ;
        RECT 287.765 101.780 287.975 102.430 ;
        RECT 288.715 102.310 288.885 102.900 ;
        RECT 290.105 102.730 290.275 103.110 ;
        RECT 291.210 102.990 291.380 103.450 ;
        RECT 291.550 103.160 291.920 103.620 ;
        RECT 292.215 103.020 292.385 103.360 ;
        RECT 292.555 103.190 292.885 103.620 ;
        RECT 293.120 103.020 293.290 103.360 ;
        RECT 289.055 102.560 290.275 102.730 ;
        RECT 290.445 102.650 290.905 102.940 ;
        RECT 291.210 102.820 291.770 102.990 ;
        RECT 292.215 102.850 293.290 103.020 ;
        RECT 293.460 103.120 294.140 103.450 ;
        RECT 294.355 103.120 294.605 103.450 ;
        RECT 294.775 103.160 295.025 103.620 ;
        RECT 291.600 102.680 291.770 102.820 ;
        RECT 290.445 102.640 291.410 102.650 ;
        RECT 290.105 102.470 290.275 102.560 ;
        RECT 290.735 102.480 291.410 102.640 ;
        RECT 288.145 102.280 288.885 102.310 ;
        RECT 288.145 101.980 289.060 102.280 ;
        RECT 288.735 101.805 289.060 101.980 ;
        RECT 287.765 101.250 288.020 101.780 ;
        RECT 288.190 101.070 288.495 101.530 ;
        RECT 288.740 101.450 289.060 101.805 ;
        RECT 289.230 102.020 289.770 102.390 ;
        RECT 290.105 102.300 290.510 102.470 ;
        RECT 289.230 101.620 289.470 102.020 ;
        RECT 289.950 101.850 290.170 102.130 ;
        RECT 289.640 101.680 290.170 101.850 ;
        RECT 289.640 101.450 289.810 101.680 ;
        RECT 290.340 101.520 290.510 102.300 ;
        RECT 290.680 101.690 291.030 102.310 ;
        RECT 291.200 101.690 291.410 102.480 ;
        RECT 291.600 102.510 293.100 102.680 ;
        RECT 291.600 101.820 291.770 102.510 ;
        RECT 293.460 102.340 293.630 103.120 ;
        RECT 294.435 102.990 294.605 103.120 ;
        RECT 291.940 102.170 293.630 102.340 ;
        RECT 293.800 102.560 294.265 102.950 ;
        RECT 294.435 102.820 294.830 102.990 ;
        RECT 291.940 101.990 292.110 102.170 ;
        RECT 288.740 101.280 289.810 101.450 ;
        RECT 289.980 101.070 290.170 101.510 ;
        RECT 290.340 101.240 291.290 101.520 ;
        RECT 291.600 101.430 291.860 101.820 ;
        RECT 292.280 101.750 293.070 102.000 ;
        RECT 291.510 101.260 291.860 101.430 ;
        RECT 292.070 101.070 292.400 101.530 ;
        RECT 293.275 101.460 293.445 102.170 ;
        RECT 293.800 101.970 293.970 102.560 ;
        RECT 293.615 101.750 293.970 101.970 ;
        RECT 294.140 101.750 294.490 102.370 ;
        RECT 294.660 101.460 294.830 102.820 ;
        RECT 295.195 102.650 295.520 103.435 ;
        RECT 295.000 101.600 295.460 102.650 ;
        RECT 293.275 101.290 294.130 101.460 ;
        RECT 294.335 101.290 294.830 101.460 ;
        RECT 295.000 101.070 295.330 101.430 ;
        RECT 295.690 101.330 295.860 103.450 ;
        RECT 296.030 103.120 296.360 103.620 ;
        RECT 296.530 102.950 296.785 103.450 ;
        RECT 296.035 102.780 296.785 102.950 ;
        RECT 296.035 101.790 296.265 102.780 ;
        RECT 296.435 101.960 296.785 102.610 ;
        RECT 296.965 102.480 297.300 103.450 ;
        RECT 297.470 102.480 297.640 103.620 ;
        RECT 297.810 103.280 299.840 103.450 ;
        RECT 296.965 101.810 297.135 102.480 ;
        RECT 297.810 102.310 297.980 103.280 ;
        RECT 297.305 101.980 297.560 102.310 ;
        RECT 297.785 101.980 297.980 102.310 ;
        RECT 298.150 102.940 299.275 103.110 ;
        RECT 297.390 101.810 297.560 101.980 ;
        RECT 298.150 101.810 298.320 102.940 ;
        RECT 296.035 101.620 296.785 101.790 ;
        RECT 296.030 101.070 296.360 101.450 ;
        RECT 296.530 101.330 296.785 101.620 ;
        RECT 296.965 101.240 297.220 101.810 ;
        RECT 297.390 101.640 298.320 101.810 ;
        RECT 298.490 102.600 299.500 102.770 ;
        RECT 298.490 101.800 298.660 102.600 ;
        RECT 298.145 101.605 298.320 101.640 ;
        RECT 297.390 101.070 297.720 101.470 ;
        RECT 298.145 101.240 298.675 101.605 ;
        RECT 298.865 101.580 299.140 102.400 ;
        RECT 298.860 101.410 299.140 101.580 ;
        RECT 298.865 101.240 299.140 101.410 ;
        RECT 299.310 101.240 299.500 102.600 ;
        RECT 299.670 102.615 299.840 103.280 ;
        RECT 300.010 102.860 300.180 103.620 ;
        RECT 300.415 102.860 300.930 103.270 ;
        RECT 299.670 102.425 300.420 102.615 ;
        RECT 300.590 102.050 300.930 102.860 ;
        RECT 301.105 102.470 301.365 103.620 ;
        RECT 301.540 102.545 301.795 103.450 ;
        RECT 301.965 102.860 302.295 103.620 ;
        RECT 302.510 102.690 302.680 103.450 ;
        RECT 299.700 101.880 300.930 102.050 ;
        RECT 299.680 101.070 300.190 101.605 ;
        RECT 300.410 101.275 300.655 101.880 ;
        RECT 301.105 101.070 301.365 101.910 ;
        RECT 301.540 101.815 301.710 102.545 ;
        RECT 301.965 102.520 302.680 102.690 ;
        RECT 301.965 102.310 302.135 102.520 ;
        RECT 303.860 102.455 304.150 103.620 ;
        RECT 304.325 102.480 304.660 103.450 ;
        RECT 304.830 102.480 305.000 103.620 ;
        RECT 305.170 103.280 307.200 103.450 ;
        RECT 301.880 101.980 302.135 102.310 ;
        RECT 301.540 101.240 301.795 101.815 ;
        RECT 301.965 101.790 302.135 101.980 ;
        RECT 302.415 101.970 302.770 102.340 ;
        RECT 304.325 101.810 304.495 102.480 ;
        RECT 305.170 102.310 305.340 103.280 ;
        RECT 304.665 101.980 304.920 102.310 ;
        RECT 305.145 101.980 305.340 102.310 ;
        RECT 305.510 102.940 306.635 103.110 ;
        RECT 304.750 101.810 304.920 101.980 ;
        RECT 305.510 101.810 305.680 102.940 ;
        RECT 301.965 101.620 302.680 101.790 ;
        RECT 301.965 101.070 302.295 101.450 ;
        RECT 302.510 101.240 302.680 101.620 ;
        RECT 303.860 101.070 304.150 101.795 ;
        RECT 304.325 101.240 304.580 101.810 ;
        RECT 304.750 101.640 305.680 101.810 ;
        RECT 305.850 102.600 306.860 102.770 ;
        RECT 305.850 101.800 306.020 102.600 ;
        RECT 306.225 102.260 306.500 102.400 ;
        RECT 306.220 102.090 306.500 102.260 ;
        RECT 305.505 101.605 305.680 101.640 ;
        RECT 304.750 101.070 305.080 101.470 ;
        RECT 305.505 101.240 306.035 101.605 ;
        RECT 306.225 101.240 306.500 102.090 ;
        RECT 306.670 101.240 306.860 102.600 ;
        RECT 307.030 102.615 307.200 103.280 ;
        RECT 307.370 102.860 307.540 103.620 ;
        RECT 307.775 102.860 308.290 103.270 ;
        RECT 307.030 102.425 307.780 102.615 ;
        RECT 307.950 102.050 308.290 102.860 ;
        RECT 308.460 102.530 309.670 103.620 ;
        RECT 307.060 101.880 308.290 102.050 ;
        RECT 307.040 101.070 307.550 101.605 ;
        RECT 307.770 101.275 308.015 101.880 ;
        RECT 308.460 101.820 308.980 102.360 ;
        RECT 309.150 101.990 309.670 102.530 ;
        RECT 309.840 102.530 311.050 103.620 ;
        RECT 309.840 101.990 310.360 102.530 ;
        RECT 310.530 101.820 311.050 102.360 ;
        RECT 308.460 101.070 309.670 101.820 ;
        RECT 309.840 101.070 311.050 101.820 ;
        RECT 162.095 100.900 311.135 101.070 ;
        RECT 162.180 100.150 163.390 100.900 ;
        RECT 162.180 99.610 162.700 100.150 ;
        RECT 164.485 100.060 164.745 100.900 ;
        RECT 164.920 100.155 165.175 100.730 ;
        RECT 165.345 100.520 165.675 100.900 ;
        RECT 165.890 100.350 166.060 100.730 ;
        RECT 165.345 100.180 166.060 100.350 ;
        RECT 167.245 100.350 167.500 100.640 ;
        RECT 167.670 100.520 168.000 100.900 ;
        RECT 167.245 100.180 167.995 100.350 ;
        RECT 162.870 99.440 163.390 99.980 ;
        RECT 162.180 98.350 163.390 99.440 ;
        RECT 164.485 98.350 164.745 99.500 ;
        RECT 164.920 99.425 165.090 100.155 ;
        RECT 165.345 99.990 165.515 100.180 ;
        RECT 165.260 99.660 165.515 99.990 ;
        RECT 165.345 99.450 165.515 99.660 ;
        RECT 165.795 99.630 166.150 100.000 ;
        RECT 164.920 98.520 165.175 99.425 ;
        RECT 165.345 99.280 166.060 99.450 ;
        RECT 167.245 99.360 167.595 100.010 ;
        RECT 165.345 98.350 165.675 99.110 ;
        RECT 165.890 98.520 166.060 99.280 ;
        RECT 167.765 99.190 167.995 100.180 ;
        RECT 167.245 99.020 167.995 99.190 ;
        RECT 167.245 98.520 167.500 99.020 ;
        RECT 167.670 98.350 168.000 98.850 ;
        RECT 168.170 98.520 168.340 100.640 ;
        RECT 168.700 100.540 169.030 100.900 ;
        RECT 169.200 100.510 169.695 100.680 ;
        RECT 169.900 100.510 170.755 100.680 ;
        RECT 168.570 99.320 169.030 100.370 ;
        RECT 168.510 98.535 168.835 99.320 ;
        RECT 169.200 99.150 169.370 100.510 ;
        RECT 169.540 99.600 169.890 100.220 ;
        RECT 170.060 100.000 170.415 100.220 ;
        RECT 170.060 99.410 170.230 100.000 ;
        RECT 170.585 99.800 170.755 100.510 ;
        RECT 171.630 100.440 171.960 100.900 ;
        RECT 172.170 100.540 172.520 100.710 ;
        RECT 170.960 99.970 171.750 100.220 ;
        RECT 172.170 100.150 172.430 100.540 ;
        RECT 172.740 100.450 173.690 100.730 ;
        RECT 173.860 100.460 174.050 100.900 ;
        RECT 174.220 100.520 175.290 100.690 ;
        RECT 171.920 99.800 172.090 99.980 ;
        RECT 169.200 98.980 169.595 99.150 ;
        RECT 169.765 99.020 170.230 99.410 ;
        RECT 170.400 99.630 172.090 99.800 ;
        RECT 169.425 98.850 169.595 98.980 ;
        RECT 170.400 98.850 170.570 99.630 ;
        RECT 172.260 99.460 172.430 100.150 ;
        RECT 170.930 99.290 172.430 99.460 ;
        RECT 172.620 99.490 172.830 100.280 ;
        RECT 173.000 99.660 173.350 100.280 ;
        RECT 173.520 99.670 173.690 100.450 ;
        RECT 174.220 100.290 174.390 100.520 ;
        RECT 173.860 100.120 174.390 100.290 ;
        RECT 173.860 99.840 174.080 100.120 ;
        RECT 174.560 99.950 174.800 100.350 ;
        RECT 173.520 99.500 173.925 99.670 ;
        RECT 174.260 99.580 174.800 99.950 ;
        RECT 174.970 100.165 175.290 100.520 ;
        RECT 175.535 100.440 175.840 100.900 ;
        RECT 176.010 100.190 176.260 100.720 ;
        RECT 174.970 99.990 175.295 100.165 ;
        RECT 174.970 99.690 175.885 99.990 ;
        RECT 175.145 99.660 175.885 99.690 ;
        RECT 172.620 99.330 173.295 99.490 ;
        RECT 173.755 99.410 173.925 99.500 ;
        RECT 172.620 99.320 173.585 99.330 ;
        RECT 172.260 99.150 172.430 99.290 ;
        RECT 169.005 98.350 169.255 98.810 ;
        RECT 169.425 98.520 169.675 98.850 ;
        RECT 169.890 98.520 170.570 98.850 ;
        RECT 170.740 98.950 171.815 99.120 ;
        RECT 172.260 98.980 172.820 99.150 ;
        RECT 173.125 99.030 173.585 99.320 ;
        RECT 173.755 99.240 174.975 99.410 ;
        RECT 170.740 98.610 170.910 98.950 ;
        RECT 171.145 98.350 171.475 98.780 ;
        RECT 171.645 98.610 171.815 98.950 ;
        RECT 172.110 98.350 172.480 98.810 ;
        RECT 172.650 98.520 172.820 98.980 ;
        RECT 173.755 98.860 173.925 99.240 ;
        RECT 175.145 99.070 175.315 99.660 ;
        RECT 176.055 99.540 176.260 100.190 ;
        RECT 176.430 100.145 176.680 100.900 ;
        RECT 176.905 100.160 177.160 100.730 ;
        RECT 177.330 100.500 177.660 100.900 ;
        RECT 178.085 100.365 178.615 100.730 ;
        RECT 178.085 100.330 178.260 100.365 ;
        RECT 177.330 100.160 178.260 100.330 ;
        RECT 173.055 98.520 173.925 98.860 ;
        RECT 174.515 98.900 175.315 99.070 ;
        RECT 174.095 98.350 174.345 98.810 ;
        RECT 174.515 98.610 174.685 98.900 ;
        RECT 174.865 98.350 175.195 98.730 ;
        RECT 175.535 98.350 175.840 99.490 ;
        RECT 176.010 98.660 176.260 99.540 ;
        RECT 176.905 99.490 177.075 100.160 ;
        RECT 177.330 99.990 177.500 100.160 ;
        RECT 177.245 99.660 177.500 99.990 ;
        RECT 177.725 99.660 177.920 99.990 ;
        RECT 176.430 98.350 176.680 99.490 ;
        RECT 176.905 98.520 177.240 99.490 ;
        RECT 177.410 98.350 177.580 99.490 ;
        RECT 177.750 98.690 177.920 99.660 ;
        RECT 178.090 99.030 178.260 100.160 ;
        RECT 178.430 99.370 178.600 100.170 ;
        RECT 178.805 99.880 179.080 100.730 ;
        RECT 178.800 99.710 179.080 99.880 ;
        RECT 178.805 99.570 179.080 99.710 ;
        RECT 179.250 99.370 179.440 100.730 ;
        RECT 179.620 100.365 180.130 100.900 ;
        RECT 180.350 100.090 180.595 100.695 ;
        RECT 179.640 99.920 180.870 100.090 ;
        RECT 181.965 100.060 182.225 100.900 ;
        RECT 182.400 100.155 182.655 100.730 ;
        RECT 182.825 100.520 183.155 100.900 ;
        RECT 183.370 100.350 183.540 100.730 ;
        RECT 182.825 100.180 183.540 100.350 ;
        RECT 178.430 99.200 179.440 99.370 ;
        RECT 179.610 99.355 180.360 99.545 ;
        RECT 178.090 98.860 179.215 99.030 ;
        RECT 179.610 98.690 179.780 99.355 ;
        RECT 180.530 99.110 180.870 99.920 ;
        RECT 177.750 98.520 179.780 98.690 ;
        RECT 179.950 98.350 180.120 99.110 ;
        RECT 180.355 98.700 180.870 99.110 ;
        RECT 181.965 98.350 182.225 99.500 ;
        RECT 182.400 99.425 182.570 100.155 ;
        RECT 182.825 99.990 182.995 100.180 ;
        RECT 184.075 100.090 184.320 100.695 ;
        RECT 184.540 100.365 185.050 100.900 ;
        RECT 182.740 99.660 182.995 99.990 ;
        RECT 182.825 99.450 182.995 99.660 ;
        RECT 183.275 99.630 183.630 100.000 ;
        RECT 183.800 99.920 185.030 100.090 ;
        RECT 182.400 98.520 182.655 99.425 ;
        RECT 182.825 99.280 183.540 99.450 ;
        RECT 182.825 98.350 183.155 99.110 ;
        RECT 183.370 98.520 183.540 99.280 ;
        RECT 183.800 99.110 184.140 99.920 ;
        RECT 184.310 99.355 185.060 99.545 ;
        RECT 183.800 98.700 184.315 99.110 ;
        RECT 184.550 98.350 184.720 99.110 ;
        RECT 184.890 98.690 185.060 99.355 ;
        RECT 185.230 99.370 185.420 100.730 ;
        RECT 185.590 100.560 185.865 100.730 ;
        RECT 185.590 100.390 185.870 100.560 ;
        RECT 185.590 99.570 185.865 100.390 ;
        RECT 186.055 100.365 186.585 100.730 ;
        RECT 187.010 100.500 187.340 100.900 ;
        RECT 186.410 100.330 186.585 100.365 ;
        RECT 186.070 99.370 186.240 100.170 ;
        RECT 185.230 99.200 186.240 99.370 ;
        RECT 186.410 100.160 187.340 100.330 ;
        RECT 187.510 100.160 187.765 100.730 ;
        RECT 187.940 100.175 188.230 100.900 ;
        RECT 188.405 100.350 188.660 100.640 ;
        RECT 188.830 100.520 189.160 100.900 ;
        RECT 188.405 100.180 189.155 100.350 ;
        RECT 186.410 99.030 186.580 100.160 ;
        RECT 187.170 99.990 187.340 100.160 ;
        RECT 185.455 98.860 186.580 99.030 ;
        RECT 186.750 99.660 186.945 99.990 ;
        RECT 187.170 99.660 187.425 99.990 ;
        RECT 186.750 98.690 186.920 99.660 ;
        RECT 187.595 99.490 187.765 100.160 ;
        RECT 184.890 98.520 186.920 98.690 ;
        RECT 187.090 98.350 187.260 99.490 ;
        RECT 187.430 98.520 187.765 99.490 ;
        RECT 187.940 98.350 188.230 99.515 ;
        RECT 188.405 99.360 188.755 100.010 ;
        RECT 188.925 99.190 189.155 100.180 ;
        RECT 188.405 99.020 189.155 99.190 ;
        RECT 188.405 98.520 188.660 99.020 ;
        RECT 188.830 98.350 189.160 98.850 ;
        RECT 189.330 98.520 189.500 100.640 ;
        RECT 189.860 100.540 190.190 100.900 ;
        RECT 190.360 100.510 190.855 100.680 ;
        RECT 191.060 100.510 191.915 100.680 ;
        RECT 189.730 99.320 190.190 100.370 ;
        RECT 189.670 98.535 189.995 99.320 ;
        RECT 190.360 99.150 190.530 100.510 ;
        RECT 190.700 99.600 191.050 100.220 ;
        RECT 191.220 100.000 191.575 100.220 ;
        RECT 191.220 99.410 191.390 100.000 ;
        RECT 191.745 99.800 191.915 100.510 ;
        RECT 192.790 100.440 193.120 100.900 ;
        RECT 193.330 100.540 193.680 100.710 ;
        RECT 192.120 99.970 192.910 100.220 ;
        RECT 193.330 100.150 193.590 100.540 ;
        RECT 193.900 100.450 194.850 100.730 ;
        RECT 195.020 100.460 195.210 100.900 ;
        RECT 195.380 100.520 196.450 100.690 ;
        RECT 193.080 99.800 193.250 99.980 ;
        RECT 190.360 98.980 190.755 99.150 ;
        RECT 190.925 99.020 191.390 99.410 ;
        RECT 191.560 99.630 193.250 99.800 ;
        RECT 190.585 98.850 190.755 98.980 ;
        RECT 191.560 98.850 191.730 99.630 ;
        RECT 193.420 99.460 193.590 100.150 ;
        RECT 192.090 99.290 193.590 99.460 ;
        RECT 193.780 99.490 193.990 100.280 ;
        RECT 194.160 99.660 194.510 100.280 ;
        RECT 194.680 99.670 194.850 100.450 ;
        RECT 195.380 100.290 195.550 100.520 ;
        RECT 195.020 100.120 195.550 100.290 ;
        RECT 195.020 99.840 195.240 100.120 ;
        RECT 195.720 99.950 195.960 100.350 ;
        RECT 194.680 99.500 195.085 99.670 ;
        RECT 195.420 99.580 195.960 99.950 ;
        RECT 196.130 100.165 196.450 100.520 ;
        RECT 196.695 100.440 197.000 100.900 ;
        RECT 197.170 100.190 197.425 100.720 ;
        RECT 196.130 99.990 196.455 100.165 ;
        RECT 196.130 99.690 197.045 99.990 ;
        RECT 196.305 99.660 197.045 99.690 ;
        RECT 193.780 99.330 194.455 99.490 ;
        RECT 194.915 99.410 195.085 99.500 ;
        RECT 193.780 99.320 194.745 99.330 ;
        RECT 193.420 99.150 193.590 99.290 ;
        RECT 190.165 98.350 190.415 98.810 ;
        RECT 190.585 98.520 190.835 98.850 ;
        RECT 191.050 98.520 191.730 98.850 ;
        RECT 191.900 98.950 192.975 99.120 ;
        RECT 193.420 98.980 193.980 99.150 ;
        RECT 194.285 99.030 194.745 99.320 ;
        RECT 194.915 99.240 196.135 99.410 ;
        RECT 191.900 98.610 192.070 98.950 ;
        RECT 192.305 98.350 192.635 98.780 ;
        RECT 192.805 98.610 192.975 98.950 ;
        RECT 193.270 98.350 193.640 98.810 ;
        RECT 193.810 98.520 193.980 98.980 ;
        RECT 194.915 98.860 195.085 99.240 ;
        RECT 196.305 99.070 196.475 99.660 ;
        RECT 197.215 99.540 197.425 100.190 ;
        RECT 194.215 98.520 195.085 98.860 ;
        RECT 195.675 98.900 196.475 99.070 ;
        RECT 195.255 98.350 195.505 98.810 ;
        RECT 195.675 98.610 195.845 98.900 ;
        RECT 196.025 98.350 196.355 98.730 ;
        RECT 196.695 98.350 197.000 99.490 ;
        RECT 197.170 98.660 197.425 99.540 ;
        RECT 197.605 100.160 197.860 100.730 ;
        RECT 198.030 100.500 198.360 100.900 ;
        RECT 198.785 100.365 199.315 100.730 ;
        RECT 198.785 100.330 198.960 100.365 ;
        RECT 198.030 100.160 198.960 100.330 ;
        RECT 197.605 99.490 197.775 100.160 ;
        RECT 198.030 99.990 198.200 100.160 ;
        RECT 197.945 99.660 198.200 99.990 ;
        RECT 198.425 99.660 198.620 99.990 ;
        RECT 197.605 98.520 197.940 99.490 ;
        RECT 198.110 98.350 198.280 99.490 ;
        RECT 198.450 98.690 198.620 99.660 ;
        RECT 198.790 99.030 198.960 100.160 ;
        RECT 199.130 99.370 199.300 100.170 ;
        RECT 199.505 99.880 199.780 100.730 ;
        RECT 199.500 99.710 199.780 99.880 ;
        RECT 199.505 99.570 199.780 99.710 ;
        RECT 199.950 99.370 200.140 100.730 ;
        RECT 200.320 100.365 200.830 100.900 ;
        RECT 201.050 100.090 201.295 100.695 ;
        RECT 201.740 100.150 202.950 100.900 ;
        RECT 203.125 100.190 203.380 100.720 ;
        RECT 203.550 100.440 203.855 100.900 ;
        RECT 204.100 100.520 205.170 100.690 ;
        RECT 200.340 99.920 201.570 100.090 ;
        RECT 199.130 99.200 200.140 99.370 ;
        RECT 200.310 99.355 201.060 99.545 ;
        RECT 198.790 98.860 199.915 99.030 ;
        RECT 200.310 98.690 200.480 99.355 ;
        RECT 201.230 99.110 201.570 99.920 ;
        RECT 201.740 99.610 202.260 100.150 ;
        RECT 202.430 99.440 202.950 99.980 ;
        RECT 198.450 98.520 200.480 98.690 ;
        RECT 200.650 98.350 200.820 99.110 ;
        RECT 201.055 98.700 201.570 99.110 ;
        RECT 201.740 98.350 202.950 99.440 ;
        RECT 203.125 99.540 203.335 100.190 ;
        RECT 204.100 100.165 204.420 100.520 ;
        RECT 204.095 99.990 204.420 100.165 ;
        RECT 203.505 99.690 204.420 99.990 ;
        RECT 204.590 99.950 204.830 100.350 ;
        RECT 205.000 100.290 205.170 100.520 ;
        RECT 205.340 100.460 205.530 100.900 ;
        RECT 205.700 100.450 206.650 100.730 ;
        RECT 206.870 100.540 207.220 100.710 ;
        RECT 205.000 100.120 205.530 100.290 ;
        RECT 203.505 99.660 204.245 99.690 ;
        RECT 203.125 98.660 203.380 99.540 ;
        RECT 203.550 98.350 203.855 99.490 ;
        RECT 204.075 99.070 204.245 99.660 ;
        RECT 204.590 99.580 205.130 99.950 ;
        RECT 205.310 99.840 205.530 100.120 ;
        RECT 205.700 99.670 205.870 100.450 ;
        RECT 205.465 99.500 205.870 99.670 ;
        RECT 206.040 99.660 206.390 100.280 ;
        RECT 205.465 99.410 205.635 99.500 ;
        RECT 206.560 99.490 206.770 100.280 ;
        RECT 204.415 99.240 205.635 99.410 ;
        RECT 206.095 99.330 206.770 99.490 ;
        RECT 204.075 98.900 204.875 99.070 ;
        RECT 204.195 98.350 204.525 98.730 ;
        RECT 204.705 98.610 204.875 98.900 ;
        RECT 205.465 98.860 205.635 99.240 ;
        RECT 205.805 99.320 206.770 99.330 ;
        RECT 206.960 100.150 207.220 100.540 ;
        RECT 207.430 100.440 207.760 100.900 ;
        RECT 208.635 100.510 209.490 100.680 ;
        RECT 209.695 100.510 210.190 100.680 ;
        RECT 210.360 100.540 210.690 100.900 ;
        RECT 206.960 99.460 207.130 100.150 ;
        RECT 207.300 99.800 207.470 99.980 ;
        RECT 207.640 99.970 208.430 100.220 ;
        RECT 208.635 99.800 208.805 100.510 ;
        RECT 208.975 100.000 209.330 100.220 ;
        RECT 207.300 99.630 208.990 99.800 ;
        RECT 205.805 99.030 206.265 99.320 ;
        RECT 206.960 99.290 208.460 99.460 ;
        RECT 206.960 99.150 207.130 99.290 ;
        RECT 206.570 98.980 207.130 99.150 ;
        RECT 205.045 98.350 205.295 98.810 ;
        RECT 205.465 98.520 206.335 98.860 ;
        RECT 206.570 98.520 206.740 98.980 ;
        RECT 207.575 98.950 208.650 99.120 ;
        RECT 206.910 98.350 207.280 98.810 ;
        RECT 207.575 98.610 207.745 98.950 ;
        RECT 207.915 98.350 208.245 98.780 ;
        RECT 208.480 98.610 208.650 98.950 ;
        RECT 208.820 98.850 208.990 99.630 ;
        RECT 209.160 99.410 209.330 100.000 ;
        RECT 209.500 99.600 209.850 100.220 ;
        RECT 209.160 99.020 209.625 99.410 ;
        RECT 210.020 99.150 210.190 100.510 ;
        RECT 210.360 99.320 210.820 100.370 ;
        RECT 209.795 98.980 210.190 99.150 ;
        RECT 209.795 98.850 209.965 98.980 ;
        RECT 208.820 98.520 209.500 98.850 ;
        RECT 209.715 98.520 209.965 98.850 ;
        RECT 210.135 98.350 210.385 98.810 ;
        RECT 210.555 98.535 210.880 99.320 ;
        RECT 211.050 98.520 211.220 100.640 ;
        RECT 211.390 100.520 211.720 100.900 ;
        RECT 211.890 100.350 212.145 100.640 ;
        RECT 211.395 100.180 212.145 100.350 ;
        RECT 211.395 99.190 211.625 100.180 ;
        RECT 212.320 100.150 213.530 100.900 ;
        RECT 213.700 100.175 213.990 100.900 ;
        RECT 211.795 99.360 212.145 100.010 ;
        RECT 212.320 99.610 212.840 100.150 ;
        RECT 214.165 100.060 214.425 100.900 ;
        RECT 214.600 100.155 214.855 100.730 ;
        RECT 215.025 100.520 215.355 100.900 ;
        RECT 215.570 100.350 215.740 100.730 ;
        RECT 215.025 100.180 215.740 100.350 ;
        RECT 213.010 99.440 213.530 99.980 ;
        RECT 211.395 99.020 212.145 99.190 ;
        RECT 211.390 98.350 211.720 98.850 ;
        RECT 211.890 98.520 212.145 99.020 ;
        RECT 212.320 98.350 213.530 99.440 ;
        RECT 213.700 98.350 213.990 99.515 ;
        RECT 214.165 98.350 214.425 99.500 ;
        RECT 214.600 99.425 214.770 100.155 ;
        RECT 215.025 99.990 215.195 100.180 ;
        RECT 216.000 100.130 217.670 100.900 ;
        RECT 217.845 100.350 218.100 100.640 ;
        RECT 218.270 100.520 218.600 100.900 ;
        RECT 217.845 100.180 218.595 100.350 ;
        RECT 214.940 99.660 215.195 99.990 ;
        RECT 215.025 99.450 215.195 99.660 ;
        RECT 215.475 99.630 215.830 100.000 ;
        RECT 216.000 99.610 216.750 100.130 ;
        RECT 214.600 98.520 214.855 99.425 ;
        RECT 215.025 99.280 215.740 99.450 ;
        RECT 216.920 99.440 217.670 99.960 ;
        RECT 215.025 98.350 215.355 99.110 ;
        RECT 215.570 98.520 215.740 99.280 ;
        RECT 216.000 98.350 217.670 99.440 ;
        RECT 217.845 99.360 218.195 100.010 ;
        RECT 218.365 99.190 218.595 100.180 ;
        RECT 217.845 99.020 218.595 99.190 ;
        RECT 217.845 98.520 218.100 99.020 ;
        RECT 218.270 98.350 218.600 98.850 ;
        RECT 218.770 98.520 218.940 100.640 ;
        RECT 219.300 100.540 219.630 100.900 ;
        RECT 219.800 100.510 220.295 100.680 ;
        RECT 220.500 100.510 221.355 100.680 ;
        RECT 219.170 99.320 219.630 100.370 ;
        RECT 219.110 98.535 219.435 99.320 ;
        RECT 219.800 99.150 219.970 100.510 ;
        RECT 220.140 99.600 220.490 100.220 ;
        RECT 220.660 100.000 221.015 100.220 ;
        RECT 220.660 99.410 220.830 100.000 ;
        RECT 221.185 99.800 221.355 100.510 ;
        RECT 222.230 100.440 222.560 100.900 ;
        RECT 222.770 100.540 223.120 100.710 ;
        RECT 221.560 99.970 222.350 100.220 ;
        RECT 222.770 100.150 223.030 100.540 ;
        RECT 223.340 100.450 224.290 100.730 ;
        RECT 224.460 100.460 224.650 100.900 ;
        RECT 224.820 100.520 225.890 100.690 ;
        RECT 222.520 99.800 222.690 99.980 ;
        RECT 219.800 98.980 220.195 99.150 ;
        RECT 220.365 99.020 220.830 99.410 ;
        RECT 221.000 99.630 222.690 99.800 ;
        RECT 220.025 98.850 220.195 98.980 ;
        RECT 221.000 98.850 221.170 99.630 ;
        RECT 222.860 99.460 223.030 100.150 ;
        RECT 221.530 99.290 223.030 99.460 ;
        RECT 223.220 99.490 223.430 100.280 ;
        RECT 223.600 99.660 223.950 100.280 ;
        RECT 224.120 99.670 224.290 100.450 ;
        RECT 224.820 100.290 224.990 100.520 ;
        RECT 224.460 100.120 224.990 100.290 ;
        RECT 224.460 99.840 224.680 100.120 ;
        RECT 225.160 99.950 225.400 100.350 ;
        RECT 224.120 99.500 224.525 99.670 ;
        RECT 224.860 99.580 225.400 99.950 ;
        RECT 225.570 100.165 225.890 100.520 ;
        RECT 226.135 100.440 226.440 100.900 ;
        RECT 226.610 100.190 226.865 100.720 ;
        RECT 225.570 99.990 225.895 100.165 ;
        RECT 225.570 99.690 226.485 99.990 ;
        RECT 225.745 99.660 226.485 99.690 ;
        RECT 223.220 99.330 223.895 99.490 ;
        RECT 224.355 99.410 224.525 99.500 ;
        RECT 223.220 99.320 224.185 99.330 ;
        RECT 222.860 99.150 223.030 99.290 ;
        RECT 219.605 98.350 219.855 98.810 ;
        RECT 220.025 98.520 220.275 98.850 ;
        RECT 220.490 98.520 221.170 98.850 ;
        RECT 221.340 98.950 222.415 99.120 ;
        RECT 222.860 98.980 223.420 99.150 ;
        RECT 223.725 99.030 224.185 99.320 ;
        RECT 224.355 99.240 225.575 99.410 ;
        RECT 221.340 98.610 221.510 98.950 ;
        RECT 221.745 98.350 222.075 98.780 ;
        RECT 222.245 98.610 222.415 98.950 ;
        RECT 222.710 98.350 223.080 98.810 ;
        RECT 223.250 98.520 223.420 98.980 ;
        RECT 224.355 98.860 224.525 99.240 ;
        RECT 225.745 99.070 225.915 99.660 ;
        RECT 226.655 99.540 226.865 100.190 ;
        RECT 223.655 98.520 224.525 98.860 ;
        RECT 225.115 98.900 225.915 99.070 ;
        RECT 224.695 98.350 224.945 98.810 ;
        RECT 225.115 98.610 225.285 98.900 ;
        RECT 225.465 98.350 225.795 98.730 ;
        RECT 226.135 98.350 226.440 99.490 ;
        RECT 226.610 98.660 226.865 99.540 ;
        RECT 227.040 99.955 227.380 100.730 ;
        RECT 227.550 100.440 227.720 100.900 ;
        RECT 227.960 100.465 228.320 100.730 ;
        RECT 227.960 100.460 228.315 100.465 ;
        RECT 227.960 100.450 228.310 100.460 ;
        RECT 227.960 100.445 228.305 100.450 ;
        RECT 227.960 100.435 228.300 100.445 ;
        RECT 228.950 100.440 229.120 100.900 ;
        RECT 227.960 100.430 228.295 100.435 ;
        RECT 227.960 100.420 228.285 100.430 ;
        RECT 227.960 100.410 228.275 100.420 ;
        RECT 227.960 100.270 228.260 100.410 ;
        RECT 227.550 100.080 228.260 100.270 ;
        RECT 228.450 100.270 228.780 100.350 ;
        RECT 229.290 100.270 229.630 100.730 ;
        RECT 229.800 100.355 235.145 100.900 ;
        RECT 228.450 100.080 229.630 100.270 ;
        RECT 227.040 98.520 227.320 99.955 ;
        RECT 227.550 99.510 227.835 100.080 ;
        RECT 228.020 99.680 228.490 99.910 ;
        RECT 228.660 99.890 228.990 99.910 ;
        RECT 228.660 99.710 229.110 99.890 ;
        RECT 229.300 99.710 229.630 99.910 ;
        RECT 227.550 99.295 228.700 99.510 ;
        RECT 227.490 98.350 228.200 99.125 ;
        RECT 228.370 98.520 228.700 99.295 ;
        RECT 228.895 98.595 229.110 99.710 ;
        RECT 229.400 99.370 229.630 99.710 ;
        RECT 231.385 99.525 231.725 100.355 ;
        RECT 235.320 100.130 238.830 100.900 ;
        RECT 239.460 100.175 239.750 100.900 ;
        RECT 239.925 100.350 240.180 100.640 ;
        RECT 240.350 100.520 240.680 100.900 ;
        RECT 239.925 100.180 240.675 100.350 ;
        RECT 229.290 98.350 229.620 99.070 ;
        RECT 233.205 98.785 233.555 100.035 ;
        RECT 235.320 99.610 236.970 100.130 ;
        RECT 237.140 99.440 238.830 99.960 ;
        RECT 229.800 98.350 235.145 98.785 ;
        RECT 235.320 98.350 238.830 99.440 ;
        RECT 239.460 98.350 239.750 99.515 ;
        RECT 239.925 99.360 240.275 100.010 ;
        RECT 240.445 99.190 240.675 100.180 ;
        RECT 239.925 99.020 240.675 99.190 ;
        RECT 239.925 98.520 240.180 99.020 ;
        RECT 240.350 98.350 240.680 98.850 ;
        RECT 240.850 98.520 241.020 100.640 ;
        RECT 241.380 100.540 241.710 100.900 ;
        RECT 241.880 100.510 242.375 100.680 ;
        RECT 242.580 100.510 243.435 100.680 ;
        RECT 241.250 99.320 241.710 100.370 ;
        RECT 241.190 98.535 241.515 99.320 ;
        RECT 241.880 99.150 242.050 100.510 ;
        RECT 242.220 99.600 242.570 100.220 ;
        RECT 242.740 100.000 243.095 100.220 ;
        RECT 242.740 99.410 242.910 100.000 ;
        RECT 243.265 99.800 243.435 100.510 ;
        RECT 244.310 100.440 244.640 100.900 ;
        RECT 244.850 100.540 245.200 100.710 ;
        RECT 243.640 99.970 244.430 100.220 ;
        RECT 244.850 100.150 245.110 100.540 ;
        RECT 245.420 100.450 246.370 100.730 ;
        RECT 246.540 100.460 246.730 100.900 ;
        RECT 246.900 100.520 247.970 100.690 ;
        RECT 244.600 99.800 244.770 99.980 ;
        RECT 241.880 98.980 242.275 99.150 ;
        RECT 242.445 99.020 242.910 99.410 ;
        RECT 243.080 99.630 244.770 99.800 ;
        RECT 242.105 98.850 242.275 98.980 ;
        RECT 243.080 98.850 243.250 99.630 ;
        RECT 244.940 99.460 245.110 100.150 ;
        RECT 243.610 99.290 245.110 99.460 ;
        RECT 245.300 99.490 245.510 100.280 ;
        RECT 245.680 99.660 246.030 100.280 ;
        RECT 246.200 99.670 246.370 100.450 ;
        RECT 246.900 100.290 247.070 100.520 ;
        RECT 246.540 100.120 247.070 100.290 ;
        RECT 246.540 99.840 246.760 100.120 ;
        RECT 247.240 99.950 247.480 100.350 ;
        RECT 246.200 99.500 246.605 99.670 ;
        RECT 246.940 99.580 247.480 99.950 ;
        RECT 247.650 100.165 247.970 100.520 ;
        RECT 248.215 100.440 248.520 100.900 ;
        RECT 248.690 100.190 248.945 100.720 ;
        RECT 247.650 99.990 247.975 100.165 ;
        RECT 247.650 99.690 248.565 99.990 ;
        RECT 247.825 99.660 248.565 99.690 ;
        RECT 245.300 99.330 245.975 99.490 ;
        RECT 246.435 99.410 246.605 99.500 ;
        RECT 245.300 99.320 246.265 99.330 ;
        RECT 244.940 99.150 245.110 99.290 ;
        RECT 241.685 98.350 241.935 98.810 ;
        RECT 242.105 98.520 242.355 98.850 ;
        RECT 242.570 98.520 243.250 98.850 ;
        RECT 243.420 98.950 244.495 99.120 ;
        RECT 244.940 98.980 245.500 99.150 ;
        RECT 245.805 99.030 246.265 99.320 ;
        RECT 246.435 99.240 247.655 99.410 ;
        RECT 243.420 98.610 243.590 98.950 ;
        RECT 243.825 98.350 244.155 98.780 ;
        RECT 244.325 98.610 244.495 98.950 ;
        RECT 244.790 98.350 245.160 98.810 ;
        RECT 245.330 98.520 245.500 98.980 ;
        RECT 246.435 98.860 246.605 99.240 ;
        RECT 247.825 99.070 247.995 99.660 ;
        RECT 248.735 99.540 248.945 100.190 ;
        RECT 249.125 100.350 249.380 100.640 ;
        RECT 249.550 100.520 249.880 100.900 ;
        RECT 249.125 100.180 249.875 100.350 ;
        RECT 245.735 98.520 246.605 98.860 ;
        RECT 247.195 98.900 247.995 99.070 ;
        RECT 246.775 98.350 247.025 98.810 ;
        RECT 247.195 98.610 247.365 98.900 ;
        RECT 247.545 98.350 247.875 98.730 ;
        RECT 248.215 98.350 248.520 99.490 ;
        RECT 248.690 98.660 248.945 99.540 ;
        RECT 249.125 99.360 249.475 100.010 ;
        RECT 249.645 99.190 249.875 100.180 ;
        RECT 249.125 99.020 249.875 99.190 ;
        RECT 249.125 98.520 249.380 99.020 ;
        RECT 249.550 98.350 249.880 98.850 ;
        RECT 250.050 98.520 250.220 100.640 ;
        RECT 250.580 100.540 250.910 100.900 ;
        RECT 251.080 100.510 251.575 100.680 ;
        RECT 251.780 100.510 252.635 100.680 ;
        RECT 250.450 99.320 250.910 100.370 ;
        RECT 250.390 98.535 250.715 99.320 ;
        RECT 251.080 99.150 251.250 100.510 ;
        RECT 251.420 99.600 251.770 100.220 ;
        RECT 251.940 100.000 252.295 100.220 ;
        RECT 251.940 99.410 252.110 100.000 ;
        RECT 252.465 99.800 252.635 100.510 ;
        RECT 253.510 100.440 253.840 100.900 ;
        RECT 254.050 100.540 254.400 100.710 ;
        RECT 252.840 99.970 253.630 100.220 ;
        RECT 254.050 100.150 254.310 100.540 ;
        RECT 254.620 100.450 255.570 100.730 ;
        RECT 255.740 100.460 255.930 100.900 ;
        RECT 256.100 100.520 257.170 100.690 ;
        RECT 253.800 99.800 253.970 99.980 ;
        RECT 251.080 98.980 251.475 99.150 ;
        RECT 251.645 99.020 252.110 99.410 ;
        RECT 252.280 99.630 253.970 99.800 ;
        RECT 251.305 98.850 251.475 98.980 ;
        RECT 252.280 98.850 252.450 99.630 ;
        RECT 254.140 99.460 254.310 100.150 ;
        RECT 252.810 99.290 254.310 99.460 ;
        RECT 254.500 99.490 254.710 100.280 ;
        RECT 254.880 99.660 255.230 100.280 ;
        RECT 255.400 99.670 255.570 100.450 ;
        RECT 256.100 100.290 256.270 100.520 ;
        RECT 255.740 100.120 256.270 100.290 ;
        RECT 255.740 99.840 255.960 100.120 ;
        RECT 256.440 99.950 256.680 100.350 ;
        RECT 255.400 99.500 255.805 99.670 ;
        RECT 256.140 99.580 256.680 99.950 ;
        RECT 256.850 100.165 257.170 100.520 ;
        RECT 257.415 100.440 257.720 100.900 ;
        RECT 257.890 100.190 258.145 100.720 ;
        RECT 256.850 99.990 257.175 100.165 ;
        RECT 256.850 99.690 257.765 99.990 ;
        RECT 257.025 99.660 257.765 99.690 ;
        RECT 254.500 99.330 255.175 99.490 ;
        RECT 255.635 99.410 255.805 99.500 ;
        RECT 254.500 99.320 255.465 99.330 ;
        RECT 254.140 99.150 254.310 99.290 ;
        RECT 250.885 98.350 251.135 98.810 ;
        RECT 251.305 98.520 251.555 98.850 ;
        RECT 251.770 98.520 252.450 98.850 ;
        RECT 252.620 98.950 253.695 99.120 ;
        RECT 254.140 98.980 254.700 99.150 ;
        RECT 255.005 99.030 255.465 99.320 ;
        RECT 255.635 99.240 256.855 99.410 ;
        RECT 252.620 98.610 252.790 98.950 ;
        RECT 253.025 98.350 253.355 98.780 ;
        RECT 253.525 98.610 253.695 98.950 ;
        RECT 253.990 98.350 254.360 98.810 ;
        RECT 254.530 98.520 254.700 98.980 ;
        RECT 255.635 98.860 255.805 99.240 ;
        RECT 257.025 99.070 257.195 99.660 ;
        RECT 257.935 99.540 258.145 100.190 ;
        RECT 258.325 100.060 258.585 100.900 ;
        RECT 258.760 100.155 259.015 100.730 ;
        RECT 259.185 100.520 259.515 100.900 ;
        RECT 259.730 100.350 259.900 100.730 ;
        RECT 259.185 100.180 259.900 100.350 ;
        RECT 254.935 98.520 255.805 98.860 ;
        RECT 256.395 98.900 257.195 99.070 ;
        RECT 255.975 98.350 256.225 98.810 ;
        RECT 256.395 98.610 256.565 98.900 ;
        RECT 256.745 98.350 257.075 98.730 ;
        RECT 257.415 98.350 257.720 99.490 ;
        RECT 257.890 98.660 258.145 99.540 ;
        RECT 258.325 98.350 258.585 99.500 ;
        RECT 258.760 99.425 258.930 100.155 ;
        RECT 259.185 99.990 259.355 100.180 ;
        RECT 260.160 100.130 262.750 100.900 ;
        RECT 259.100 99.660 259.355 99.990 ;
        RECT 259.185 99.450 259.355 99.660 ;
        RECT 259.635 99.630 259.990 100.000 ;
        RECT 260.160 99.610 261.370 100.130 ;
        RECT 263.385 100.060 263.645 100.900 ;
        RECT 263.820 100.155 264.075 100.730 ;
        RECT 264.245 100.520 264.575 100.900 ;
        RECT 264.790 100.350 264.960 100.730 ;
        RECT 264.245 100.180 264.960 100.350 ;
        RECT 258.760 98.520 259.015 99.425 ;
        RECT 259.185 99.280 259.900 99.450 ;
        RECT 261.540 99.440 262.750 99.960 ;
        RECT 259.185 98.350 259.515 99.110 ;
        RECT 259.730 98.520 259.900 99.280 ;
        RECT 260.160 98.350 262.750 99.440 ;
        RECT 263.385 98.350 263.645 99.500 ;
        RECT 263.820 99.425 263.990 100.155 ;
        RECT 264.245 99.990 264.415 100.180 ;
        RECT 265.220 100.175 265.510 100.900 ;
        RECT 265.680 100.150 266.890 100.900 ;
        RECT 267.065 100.160 267.320 100.730 ;
        RECT 267.490 100.500 267.820 100.900 ;
        RECT 268.245 100.365 268.775 100.730 ;
        RECT 268.965 100.560 269.240 100.730 ;
        RECT 268.960 100.390 269.240 100.560 ;
        RECT 268.245 100.330 268.420 100.365 ;
        RECT 267.490 100.160 268.420 100.330 ;
        RECT 264.160 99.660 264.415 99.990 ;
        RECT 264.245 99.450 264.415 99.660 ;
        RECT 264.695 99.630 265.050 100.000 ;
        RECT 265.680 99.610 266.200 100.150 ;
        RECT 263.820 98.520 264.075 99.425 ;
        RECT 264.245 99.280 264.960 99.450 ;
        RECT 264.245 98.350 264.575 99.110 ;
        RECT 264.790 98.520 264.960 99.280 ;
        RECT 265.220 98.350 265.510 99.515 ;
        RECT 266.370 99.440 266.890 99.980 ;
        RECT 265.680 98.350 266.890 99.440 ;
        RECT 267.065 99.490 267.235 100.160 ;
        RECT 267.490 99.990 267.660 100.160 ;
        RECT 267.405 99.660 267.660 99.990 ;
        RECT 267.885 99.660 268.080 99.990 ;
        RECT 267.065 98.520 267.400 99.490 ;
        RECT 267.570 98.350 267.740 99.490 ;
        RECT 267.910 98.690 268.080 99.660 ;
        RECT 268.250 99.030 268.420 100.160 ;
        RECT 268.590 99.370 268.760 100.170 ;
        RECT 268.965 99.570 269.240 100.390 ;
        RECT 269.410 99.370 269.600 100.730 ;
        RECT 269.780 100.365 270.290 100.900 ;
        RECT 270.510 100.090 270.755 100.695 ;
        RECT 271.665 100.350 271.920 100.640 ;
        RECT 272.090 100.520 272.420 100.900 ;
        RECT 271.665 100.180 272.415 100.350 ;
        RECT 269.800 99.920 271.030 100.090 ;
        RECT 268.590 99.200 269.600 99.370 ;
        RECT 269.770 99.355 270.520 99.545 ;
        RECT 268.250 98.860 269.375 99.030 ;
        RECT 269.770 98.690 269.940 99.355 ;
        RECT 270.690 99.110 271.030 99.920 ;
        RECT 271.665 99.360 272.015 100.010 ;
        RECT 272.185 99.190 272.415 100.180 ;
        RECT 267.910 98.520 269.940 98.690 ;
        RECT 270.110 98.350 270.280 99.110 ;
        RECT 270.515 98.700 271.030 99.110 ;
        RECT 271.665 99.020 272.415 99.190 ;
        RECT 271.665 98.520 271.920 99.020 ;
        RECT 272.090 98.350 272.420 98.850 ;
        RECT 272.590 98.520 272.760 100.640 ;
        RECT 273.120 100.540 273.450 100.900 ;
        RECT 273.620 100.510 274.115 100.680 ;
        RECT 274.320 100.510 275.175 100.680 ;
        RECT 272.990 99.320 273.450 100.370 ;
        RECT 272.930 98.535 273.255 99.320 ;
        RECT 273.620 99.150 273.790 100.510 ;
        RECT 273.960 99.600 274.310 100.220 ;
        RECT 274.480 100.000 274.835 100.220 ;
        RECT 274.480 99.410 274.650 100.000 ;
        RECT 275.005 99.800 275.175 100.510 ;
        RECT 276.050 100.440 276.380 100.900 ;
        RECT 276.590 100.540 276.940 100.710 ;
        RECT 275.380 99.970 276.170 100.220 ;
        RECT 276.590 100.150 276.850 100.540 ;
        RECT 277.160 100.450 278.110 100.730 ;
        RECT 278.280 100.460 278.470 100.900 ;
        RECT 278.640 100.520 279.710 100.690 ;
        RECT 276.340 99.800 276.510 99.980 ;
        RECT 273.620 98.980 274.015 99.150 ;
        RECT 274.185 99.020 274.650 99.410 ;
        RECT 274.820 99.630 276.510 99.800 ;
        RECT 273.845 98.850 274.015 98.980 ;
        RECT 274.820 98.850 274.990 99.630 ;
        RECT 276.680 99.460 276.850 100.150 ;
        RECT 275.350 99.290 276.850 99.460 ;
        RECT 277.040 99.490 277.250 100.280 ;
        RECT 277.420 99.660 277.770 100.280 ;
        RECT 277.940 99.670 278.110 100.450 ;
        RECT 278.640 100.290 278.810 100.520 ;
        RECT 278.280 100.120 278.810 100.290 ;
        RECT 278.280 99.840 278.500 100.120 ;
        RECT 278.980 99.950 279.220 100.350 ;
        RECT 277.940 99.500 278.345 99.670 ;
        RECT 278.680 99.580 279.220 99.950 ;
        RECT 279.390 100.165 279.710 100.520 ;
        RECT 279.955 100.440 280.260 100.900 ;
        RECT 280.430 100.190 280.685 100.720 ;
        RECT 279.390 99.990 279.715 100.165 ;
        RECT 279.390 99.690 280.305 99.990 ;
        RECT 279.565 99.660 280.305 99.690 ;
        RECT 277.040 99.330 277.715 99.490 ;
        RECT 278.175 99.410 278.345 99.500 ;
        RECT 277.040 99.320 278.005 99.330 ;
        RECT 276.680 99.150 276.850 99.290 ;
        RECT 273.425 98.350 273.675 98.810 ;
        RECT 273.845 98.520 274.095 98.850 ;
        RECT 274.310 98.520 274.990 98.850 ;
        RECT 275.160 98.950 276.235 99.120 ;
        RECT 276.680 98.980 277.240 99.150 ;
        RECT 277.545 99.030 278.005 99.320 ;
        RECT 278.175 99.240 279.395 99.410 ;
        RECT 275.160 98.610 275.330 98.950 ;
        RECT 275.565 98.350 275.895 98.780 ;
        RECT 276.065 98.610 276.235 98.950 ;
        RECT 276.530 98.350 276.900 98.810 ;
        RECT 277.070 98.520 277.240 98.980 ;
        RECT 278.175 98.860 278.345 99.240 ;
        RECT 279.565 99.070 279.735 99.660 ;
        RECT 280.475 99.540 280.685 100.190 ;
        RECT 281.135 100.090 281.380 100.695 ;
        RECT 281.600 100.365 282.110 100.900 ;
        RECT 277.475 98.520 278.345 98.860 ;
        RECT 278.935 98.900 279.735 99.070 ;
        RECT 278.515 98.350 278.765 98.810 ;
        RECT 278.935 98.610 279.105 98.900 ;
        RECT 279.285 98.350 279.615 98.730 ;
        RECT 279.955 98.350 280.260 99.490 ;
        RECT 280.430 98.660 280.685 99.540 ;
        RECT 280.860 99.920 282.090 100.090 ;
        RECT 280.860 99.110 281.200 99.920 ;
        RECT 281.370 99.355 282.120 99.545 ;
        RECT 280.860 98.700 281.375 99.110 ;
        RECT 281.610 98.350 281.780 99.110 ;
        RECT 281.950 98.690 282.120 99.355 ;
        RECT 282.290 99.370 282.480 100.730 ;
        RECT 282.650 100.560 282.925 100.730 ;
        RECT 282.650 100.390 282.930 100.560 ;
        RECT 282.650 99.570 282.925 100.390 ;
        RECT 283.115 100.365 283.645 100.730 ;
        RECT 284.070 100.500 284.400 100.900 ;
        RECT 283.470 100.330 283.645 100.365 ;
        RECT 283.130 99.370 283.300 100.170 ;
        RECT 282.290 99.200 283.300 99.370 ;
        RECT 283.470 100.160 284.400 100.330 ;
        RECT 284.570 100.160 284.825 100.730 ;
        RECT 283.470 99.030 283.640 100.160 ;
        RECT 284.230 99.990 284.400 100.160 ;
        RECT 282.515 98.860 283.640 99.030 ;
        RECT 283.810 99.660 284.005 99.990 ;
        RECT 284.230 99.660 284.485 99.990 ;
        RECT 283.810 98.690 283.980 99.660 ;
        RECT 284.655 99.490 284.825 100.160 ;
        RECT 285.005 100.060 285.265 100.900 ;
        RECT 285.440 100.155 285.695 100.730 ;
        RECT 285.865 100.520 286.195 100.900 ;
        RECT 286.410 100.350 286.580 100.730 ;
        RECT 285.865 100.180 286.580 100.350 ;
        RECT 281.950 98.520 283.980 98.690 ;
        RECT 284.150 98.350 284.320 99.490 ;
        RECT 284.490 98.520 284.825 99.490 ;
        RECT 285.005 98.350 285.265 99.500 ;
        RECT 285.440 99.425 285.610 100.155 ;
        RECT 285.865 99.990 286.035 100.180 ;
        RECT 286.845 100.060 287.105 100.900 ;
        RECT 287.280 100.155 287.535 100.730 ;
        RECT 287.705 100.520 288.035 100.900 ;
        RECT 288.250 100.350 288.420 100.730 ;
        RECT 287.705 100.180 288.420 100.350 ;
        RECT 285.780 99.660 286.035 99.990 ;
        RECT 285.865 99.450 286.035 99.660 ;
        RECT 286.315 99.630 286.670 100.000 ;
        RECT 285.440 98.520 285.695 99.425 ;
        RECT 285.865 99.280 286.580 99.450 ;
        RECT 285.865 98.350 286.195 99.110 ;
        RECT 286.410 98.520 286.580 99.280 ;
        RECT 286.845 98.350 287.105 99.500 ;
        RECT 287.280 99.425 287.450 100.155 ;
        RECT 287.705 99.990 287.875 100.180 ;
        RECT 288.685 100.060 288.945 100.900 ;
        RECT 289.120 100.155 289.375 100.730 ;
        RECT 289.545 100.520 289.875 100.900 ;
        RECT 290.090 100.350 290.260 100.730 ;
        RECT 289.545 100.180 290.260 100.350 ;
        RECT 287.620 99.660 287.875 99.990 ;
        RECT 287.705 99.450 287.875 99.660 ;
        RECT 288.155 99.630 288.510 100.000 ;
        RECT 287.280 98.520 287.535 99.425 ;
        RECT 287.705 99.280 288.420 99.450 ;
        RECT 287.705 98.350 288.035 99.110 ;
        RECT 288.250 98.520 288.420 99.280 ;
        RECT 288.685 98.350 288.945 99.500 ;
        RECT 289.120 99.425 289.290 100.155 ;
        RECT 289.545 99.990 289.715 100.180 ;
        RECT 290.980 100.175 291.270 100.900 ;
        RECT 291.445 100.160 291.700 100.730 ;
        RECT 291.870 100.500 292.200 100.900 ;
        RECT 292.625 100.365 293.155 100.730 ;
        RECT 292.625 100.330 292.800 100.365 ;
        RECT 291.870 100.160 292.800 100.330 ;
        RECT 289.460 99.660 289.715 99.990 ;
        RECT 289.545 99.450 289.715 99.660 ;
        RECT 289.995 99.630 290.350 100.000 ;
        RECT 289.120 98.520 289.375 99.425 ;
        RECT 289.545 99.280 290.260 99.450 ;
        RECT 289.545 98.350 289.875 99.110 ;
        RECT 290.090 98.520 290.260 99.280 ;
        RECT 290.980 98.350 291.270 99.515 ;
        RECT 291.445 99.490 291.615 100.160 ;
        RECT 291.870 99.990 292.040 100.160 ;
        RECT 291.785 99.660 292.040 99.990 ;
        RECT 292.265 99.660 292.460 99.990 ;
        RECT 291.445 98.520 291.780 99.490 ;
        RECT 291.950 98.350 292.120 99.490 ;
        RECT 292.290 98.690 292.460 99.660 ;
        RECT 292.630 99.030 292.800 100.160 ;
        RECT 292.970 99.370 293.140 100.170 ;
        RECT 293.345 99.880 293.620 100.730 ;
        RECT 293.340 99.710 293.620 99.880 ;
        RECT 293.345 99.570 293.620 99.710 ;
        RECT 293.790 99.370 293.980 100.730 ;
        RECT 294.160 100.365 294.670 100.900 ;
        RECT 294.890 100.090 295.135 100.695 ;
        RECT 296.045 100.350 296.300 100.640 ;
        RECT 296.470 100.520 296.800 100.900 ;
        RECT 296.045 100.180 296.795 100.350 ;
        RECT 294.180 99.920 295.410 100.090 ;
        RECT 292.970 99.200 293.980 99.370 ;
        RECT 294.150 99.355 294.900 99.545 ;
        RECT 292.630 98.860 293.755 99.030 ;
        RECT 294.150 98.690 294.320 99.355 ;
        RECT 295.070 99.110 295.410 99.920 ;
        RECT 296.045 99.360 296.395 100.010 ;
        RECT 296.565 99.190 296.795 100.180 ;
        RECT 292.290 98.520 294.320 98.690 ;
        RECT 294.490 98.350 294.660 99.110 ;
        RECT 294.895 98.700 295.410 99.110 ;
        RECT 296.045 99.020 296.795 99.190 ;
        RECT 296.045 98.520 296.300 99.020 ;
        RECT 296.470 98.350 296.800 98.850 ;
        RECT 296.970 98.520 297.140 100.640 ;
        RECT 297.500 100.540 297.830 100.900 ;
        RECT 298.000 100.510 298.495 100.680 ;
        RECT 298.700 100.510 299.555 100.680 ;
        RECT 297.370 99.320 297.830 100.370 ;
        RECT 297.310 98.535 297.635 99.320 ;
        RECT 298.000 99.150 298.170 100.510 ;
        RECT 298.340 99.600 298.690 100.220 ;
        RECT 298.860 100.000 299.215 100.220 ;
        RECT 298.860 99.410 299.030 100.000 ;
        RECT 299.385 99.800 299.555 100.510 ;
        RECT 300.430 100.440 300.760 100.900 ;
        RECT 300.970 100.540 301.320 100.710 ;
        RECT 299.760 99.970 300.550 100.220 ;
        RECT 300.970 100.150 301.230 100.540 ;
        RECT 301.540 100.450 302.490 100.730 ;
        RECT 302.660 100.460 302.850 100.900 ;
        RECT 303.020 100.520 304.090 100.690 ;
        RECT 300.720 99.800 300.890 99.980 ;
        RECT 298.000 98.980 298.395 99.150 ;
        RECT 298.565 99.020 299.030 99.410 ;
        RECT 299.200 99.630 300.890 99.800 ;
        RECT 298.225 98.850 298.395 98.980 ;
        RECT 299.200 98.850 299.370 99.630 ;
        RECT 301.060 99.460 301.230 100.150 ;
        RECT 299.730 99.290 301.230 99.460 ;
        RECT 301.420 99.490 301.630 100.280 ;
        RECT 301.800 99.660 302.150 100.280 ;
        RECT 302.320 99.670 302.490 100.450 ;
        RECT 303.020 100.290 303.190 100.520 ;
        RECT 302.660 100.120 303.190 100.290 ;
        RECT 302.660 99.840 302.880 100.120 ;
        RECT 303.360 99.950 303.600 100.350 ;
        RECT 302.320 99.500 302.725 99.670 ;
        RECT 303.060 99.580 303.600 99.950 ;
        RECT 303.770 100.165 304.090 100.520 ;
        RECT 304.335 100.440 304.640 100.900 ;
        RECT 304.810 100.190 305.065 100.720 ;
        RECT 303.770 99.990 304.095 100.165 ;
        RECT 303.770 99.690 304.685 99.990 ;
        RECT 303.945 99.660 304.685 99.690 ;
        RECT 301.420 99.330 302.095 99.490 ;
        RECT 302.555 99.410 302.725 99.500 ;
        RECT 301.420 99.320 302.385 99.330 ;
        RECT 301.060 99.150 301.230 99.290 ;
        RECT 297.805 98.350 298.055 98.810 ;
        RECT 298.225 98.520 298.475 98.850 ;
        RECT 298.690 98.520 299.370 98.850 ;
        RECT 299.540 98.950 300.615 99.120 ;
        RECT 301.060 98.980 301.620 99.150 ;
        RECT 301.925 99.030 302.385 99.320 ;
        RECT 302.555 99.240 303.775 99.410 ;
        RECT 299.540 98.610 299.710 98.950 ;
        RECT 299.945 98.350 300.275 98.780 ;
        RECT 300.445 98.610 300.615 98.950 ;
        RECT 300.910 98.350 301.280 98.810 ;
        RECT 301.450 98.520 301.620 98.980 ;
        RECT 302.555 98.860 302.725 99.240 ;
        RECT 303.945 99.070 304.115 99.660 ;
        RECT 304.855 99.540 305.065 100.190 ;
        RECT 305.330 100.350 305.500 100.730 ;
        RECT 305.715 100.520 306.045 100.900 ;
        RECT 305.330 100.180 306.045 100.350 ;
        RECT 305.240 99.630 305.595 100.000 ;
        RECT 305.875 99.990 306.045 100.180 ;
        RECT 306.215 100.155 306.470 100.730 ;
        RECT 305.875 99.660 306.130 99.990 ;
        RECT 301.855 98.520 302.725 98.860 ;
        RECT 303.315 98.900 304.115 99.070 ;
        RECT 302.895 98.350 303.145 98.810 ;
        RECT 303.315 98.610 303.485 98.900 ;
        RECT 303.665 98.350 303.995 98.730 ;
        RECT 304.335 98.350 304.640 99.490 ;
        RECT 304.810 98.660 305.065 99.540 ;
        RECT 305.875 99.450 306.045 99.660 ;
        RECT 305.330 99.280 306.045 99.450 ;
        RECT 306.300 99.425 306.470 100.155 ;
        RECT 306.645 100.060 306.905 100.900 ;
        RECT 307.170 100.350 307.340 100.730 ;
        RECT 307.555 100.520 307.885 100.900 ;
        RECT 307.170 100.180 307.885 100.350 ;
        RECT 307.080 99.630 307.435 100.000 ;
        RECT 307.715 99.990 307.885 100.180 ;
        RECT 308.055 100.155 308.310 100.730 ;
        RECT 307.715 99.660 307.970 99.990 ;
        RECT 305.330 98.520 305.500 99.280 ;
        RECT 305.715 98.350 306.045 99.110 ;
        RECT 306.215 98.520 306.470 99.425 ;
        RECT 306.645 98.350 306.905 99.500 ;
        RECT 307.715 99.450 307.885 99.660 ;
        RECT 307.170 99.280 307.885 99.450 ;
        RECT 308.140 99.425 308.310 100.155 ;
        RECT 308.485 100.060 308.745 100.900 ;
        RECT 309.840 100.150 311.050 100.900 ;
        RECT 307.170 98.520 307.340 99.280 ;
        RECT 307.555 98.350 307.885 99.110 ;
        RECT 308.055 98.520 308.310 99.425 ;
        RECT 308.485 98.350 308.745 99.500 ;
        RECT 309.840 99.440 310.360 99.980 ;
        RECT 310.530 99.610 311.050 100.150 ;
        RECT 309.840 98.350 311.050 99.440 ;
        RECT 162.095 98.180 311.135 98.350 ;
        RECT 162.180 97.090 163.390 98.180 ;
        RECT 162.180 96.380 162.700 96.920 ;
        RECT 162.870 96.550 163.390 97.090 ;
        RECT 164.025 97.030 164.285 98.180 ;
        RECT 164.460 97.105 164.715 98.010 ;
        RECT 164.885 97.420 165.215 98.180 ;
        RECT 165.430 97.250 165.600 98.010 ;
        RECT 162.180 95.630 163.390 96.380 ;
        RECT 164.025 95.630 164.285 96.470 ;
        RECT 164.460 96.375 164.630 97.105 ;
        RECT 164.885 97.080 165.600 97.250 ;
        RECT 164.885 96.870 165.055 97.080 ;
        RECT 165.865 97.030 166.125 98.180 ;
        RECT 166.300 97.105 166.555 98.010 ;
        RECT 166.725 97.420 167.055 98.180 ;
        RECT 167.270 97.250 167.440 98.010 ;
        RECT 164.800 96.540 165.055 96.870 ;
        RECT 164.460 95.800 164.715 96.375 ;
        RECT 164.885 96.350 165.055 96.540 ;
        RECT 165.335 96.530 165.690 96.900 ;
        RECT 164.885 96.180 165.600 96.350 ;
        RECT 164.885 95.630 165.215 96.010 ;
        RECT 165.430 95.800 165.600 96.180 ;
        RECT 165.865 95.630 166.125 96.470 ;
        RECT 166.300 96.375 166.470 97.105 ;
        RECT 166.725 97.080 167.440 97.250 ;
        RECT 167.700 97.090 170.290 98.180 ;
        RECT 166.725 96.870 166.895 97.080 ;
        RECT 166.640 96.540 166.895 96.870 ;
        RECT 166.300 95.800 166.555 96.375 ;
        RECT 166.725 96.350 166.895 96.540 ;
        RECT 167.175 96.530 167.530 96.900 ;
        RECT 167.700 96.400 168.910 96.920 ;
        RECT 169.080 96.570 170.290 97.090 ;
        RECT 170.925 97.040 171.260 98.010 ;
        RECT 171.430 97.040 171.600 98.180 ;
        RECT 171.770 97.840 173.800 98.010 ;
        RECT 166.725 96.180 167.440 96.350 ;
        RECT 166.725 95.630 167.055 96.010 ;
        RECT 167.270 95.800 167.440 96.180 ;
        RECT 167.700 95.630 170.290 96.400 ;
        RECT 170.925 96.370 171.095 97.040 ;
        RECT 171.770 96.870 171.940 97.840 ;
        RECT 171.265 96.540 171.520 96.870 ;
        RECT 171.745 96.540 171.940 96.870 ;
        RECT 172.110 97.500 173.235 97.670 ;
        RECT 171.350 96.370 171.520 96.540 ;
        RECT 172.110 96.370 172.280 97.500 ;
        RECT 170.925 95.800 171.180 96.370 ;
        RECT 171.350 96.200 172.280 96.370 ;
        RECT 172.450 97.160 173.460 97.330 ;
        RECT 172.450 96.360 172.620 97.160 ;
        RECT 172.825 96.480 173.100 96.960 ;
        RECT 172.820 96.310 173.100 96.480 ;
        RECT 172.105 96.165 172.280 96.200 ;
        RECT 171.350 95.630 171.680 96.030 ;
        RECT 172.105 95.800 172.635 96.165 ;
        RECT 172.825 95.800 173.100 96.310 ;
        RECT 173.270 95.800 173.460 97.160 ;
        RECT 173.630 97.175 173.800 97.840 ;
        RECT 173.970 97.420 174.140 98.180 ;
        RECT 174.375 97.420 174.890 97.830 ;
        RECT 173.630 96.985 174.380 97.175 ;
        RECT 174.550 96.610 174.890 97.420 ;
        RECT 175.060 97.015 175.350 98.180 ;
        RECT 175.525 97.040 175.860 98.010 ;
        RECT 176.030 97.040 176.200 98.180 ;
        RECT 176.370 97.840 178.400 98.010 ;
        RECT 173.660 96.440 174.890 96.610 ;
        RECT 173.640 95.630 174.150 96.165 ;
        RECT 174.370 95.835 174.615 96.440 ;
        RECT 175.525 96.370 175.695 97.040 ;
        RECT 176.370 96.870 176.540 97.840 ;
        RECT 175.865 96.540 176.120 96.870 ;
        RECT 176.345 96.540 176.540 96.870 ;
        RECT 176.710 97.500 177.835 97.670 ;
        RECT 175.950 96.370 176.120 96.540 ;
        RECT 176.710 96.370 176.880 97.500 ;
        RECT 175.060 95.630 175.350 96.355 ;
        RECT 175.525 95.800 175.780 96.370 ;
        RECT 175.950 96.200 176.880 96.370 ;
        RECT 177.050 97.160 178.060 97.330 ;
        RECT 177.050 96.360 177.220 97.160 ;
        RECT 177.425 96.480 177.700 96.960 ;
        RECT 177.420 96.310 177.700 96.480 ;
        RECT 176.705 96.165 176.880 96.200 ;
        RECT 175.950 95.630 176.280 96.030 ;
        RECT 176.705 95.800 177.235 96.165 ;
        RECT 177.425 95.800 177.700 96.310 ;
        RECT 177.870 95.800 178.060 97.160 ;
        RECT 178.230 97.175 178.400 97.840 ;
        RECT 178.570 97.420 178.740 98.180 ;
        RECT 178.975 97.420 179.490 97.830 ;
        RECT 178.230 96.985 178.980 97.175 ;
        RECT 179.150 96.610 179.490 97.420 ;
        RECT 179.660 97.090 182.250 98.180 ;
        RECT 178.260 96.440 179.490 96.610 ;
        RECT 178.240 95.630 178.750 96.165 ;
        RECT 178.970 95.835 179.215 96.440 ;
        RECT 179.660 96.400 180.870 96.920 ;
        RECT 181.040 96.570 182.250 97.090 ;
        RECT 182.880 96.575 183.160 98.010 ;
        RECT 183.330 97.405 184.040 98.180 ;
        RECT 184.210 97.235 184.540 98.010 ;
        RECT 183.390 97.020 184.540 97.235 ;
        RECT 179.660 95.630 182.250 96.400 ;
        RECT 182.880 95.800 183.220 96.575 ;
        RECT 183.390 96.450 183.675 97.020 ;
        RECT 183.860 96.620 184.330 96.850 ;
        RECT 184.735 96.820 184.950 97.935 ;
        RECT 185.130 97.460 185.460 98.180 ;
        RECT 185.240 96.820 185.470 97.160 ;
        RECT 185.640 97.090 187.310 98.180 ;
        RECT 184.500 96.640 184.950 96.820 ;
        RECT 184.500 96.620 184.830 96.640 ;
        RECT 185.140 96.620 185.470 96.820 ;
        RECT 183.390 96.260 184.100 96.450 ;
        RECT 183.800 96.120 184.100 96.260 ;
        RECT 184.290 96.260 185.470 96.450 ;
        RECT 184.290 96.180 184.620 96.260 ;
        RECT 183.800 96.110 184.115 96.120 ;
        RECT 183.800 96.100 184.125 96.110 ;
        RECT 183.800 96.095 184.135 96.100 ;
        RECT 183.390 95.630 183.560 96.090 ;
        RECT 183.800 96.085 184.140 96.095 ;
        RECT 183.800 96.080 184.145 96.085 ;
        RECT 183.800 96.070 184.150 96.080 ;
        RECT 183.800 96.065 184.155 96.070 ;
        RECT 183.800 95.800 184.160 96.065 ;
        RECT 184.790 95.630 184.960 96.090 ;
        RECT 185.130 95.800 185.470 96.260 ;
        RECT 185.640 96.400 186.390 96.920 ;
        RECT 186.560 96.570 187.310 97.090 ;
        RECT 187.945 97.040 188.280 98.010 ;
        RECT 188.450 97.040 188.620 98.180 ;
        RECT 188.790 97.840 190.820 98.010 ;
        RECT 185.640 95.630 187.310 96.400 ;
        RECT 187.945 96.370 188.115 97.040 ;
        RECT 188.790 96.870 188.960 97.840 ;
        RECT 188.285 96.540 188.540 96.870 ;
        RECT 188.765 96.540 188.960 96.870 ;
        RECT 189.130 97.500 190.255 97.670 ;
        RECT 188.370 96.370 188.540 96.540 ;
        RECT 189.130 96.370 189.300 97.500 ;
        RECT 187.945 95.800 188.200 96.370 ;
        RECT 188.370 96.200 189.300 96.370 ;
        RECT 189.470 97.160 190.480 97.330 ;
        RECT 189.470 96.360 189.640 97.160 ;
        RECT 189.845 96.820 190.120 96.960 ;
        RECT 189.840 96.650 190.120 96.820 ;
        RECT 189.125 96.165 189.300 96.200 ;
        RECT 188.370 95.630 188.700 96.030 ;
        RECT 189.125 95.800 189.655 96.165 ;
        RECT 189.845 95.800 190.120 96.650 ;
        RECT 190.290 95.800 190.480 97.160 ;
        RECT 190.650 97.175 190.820 97.840 ;
        RECT 190.990 97.420 191.160 98.180 ;
        RECT 191.395 97.420 191.910 97.830 ;
        RECT 190.650 96.985 191.400 97.175 ;
        RECT 191.570 96.610 191.910 97.420 ;
        RECT 190.680 96.440 191.910 96.610 ;
        RECT 192.085 97.040 192.420 98.010 ;
        RECT 192.590 97.040 192.760 98.180 ;
        RECT 192.930 97.840 194.960 98.010 ;
        RECT 190.660 95.630 191.170 96.165 ;
        RECT 191.390 95.835 191.635 96.440 ;
        RECT 192.085 96.370 192.255 97.040 ;
        RECT 192.930 96.870 193.100 97.840 ;
        RECT 192.425 96.540 192.680 96.870 ;
        RECT 192.905 96.540 193.100 96.870 ;
        RECT 193.270 97.500 194.395 97.670 ;
        RECT 192.510 96.370 192.680 96.540 ;
        RECT 193.270 96.370 193.440 97.500 ;
        RECT 192.085 95.800 192.340 96.370 ;
        RECT 192.510 96.200 193.440 96.370 ;
        RECT 193.610 97.160 194.620 97.330 ;
        RECT 193.610 96.360 193.780 97.160 ;
        RECT 193.985 96.820 194.260 96.960 ;
        RECT 193.980 96.650 194.260 96.820 ;
        RECT 193.265 96.165 193.440 96.200 ;
        RECT 192.510 95.630 192.840 96.030 ;
        RECT 193.265 95.800 193.795 96.165 ;
        RECT 193.985 95.800 194.260 96.650 ;
        RECT 194.430 95.800 194.620 97.160 ;
        RECT 194.790 97.175 194.960 97.840 ;
        RECT 195.130 97.420 195.300 98.180 ;
        RECT 195.535 97.420 196.050 97.830 ;
        RECT 194.790 96.985 195.540 97.175 ;
        RECT 195.710 96.610 196.050 97.420 ;
        RECT 196.220 97.090 198.810 98.180 ;
        RECT 194.820 96.440 196.050 96.610 ;
        RECT 194.800 95.630 195.310 96.165 ;
        RECT 195.530 95.835 195.775 96.440 ;
        RECT 196.220 96.400 197.430 96.920 ;
        RECT 197.600 96.570 198.810 97.090 ;
        RECT 199.070 97.250 199.240 98.010 ;
        RECT 199.455 97.420 199.785 98.180 ;
        RECT 199.070 97.080 199.785 97.250 ;
        RECT 199.955 97.105 200.210 98.010 ;
        RECT 198.980 96.530 199.335 96.900 ;
        RECT 199.615 96.870 199.785 97.080 ;
        RECT 199.615 96.540 199.870 96.870 ;
        RECT 196.220 95.630 198.810 96.400 ;
        RECT 199.615 96.350 199.785 96.540 ;
        RECT 200.040 96.375 200.210 97.105 ;
        RECT 200.385 97.030 200.645 98.180 ;
        RECT 200.820 97.015 201.110 98.180 ;
        RECT 201.280 97.090 202.950 98.180 ;
        RECT 199.070 96.180 199.785 96.350 ;
        RECT 199.070 95.800 199.240 96.180 ;
        RECT 199.455 95.630 199.785 96.010 ;
        RECT 199.955 95.800 200.210 96.375 ;
        RECT 200.385 95.630 200.645 96.470 ;
        RECT 201.280 96.400 202.030 96.920 ;
        RECT 202.200 96.570 202.950 97.090 ;
        RECT 200.820 95.630 201.110 96.355 ;
        RECT 201.280 95.630 202.950 96.400 ;
        RECT 203.130 95.810 203.390 98.000 ;
        RECT 203.560 97.450 203.900 98.180 ;
        RECT 204.080 97.270 204.350 98.000 ;
        RECT 203.580 97.050 204.350 97.270 ;
        RECT 204.530 97.290 204.760 98.000 ;
        RECT 204.930 97.470 205.260 98.180 ;
        RECT 205.430 97.290 205.690 98.000 ;
        RECT 204.530 97.050 205.690 97.290 ;
        RECT 205.880 97.330 206.140 98.010 ;
        RECT 206.310 97.400 206.560 98.180 ;
        RECT 206.810 97.630 207.060 98.010 ;
        RECT 207.230 97.800 207.585 98.180 ;
        RECT 208.590 97.790 208.925 98.010 ;
        RECT 208.190 97.630 208.420 97.670 ;
        RECT 206.810 97.430 208.420 97.630 ;
        RECT 206.810 97.420 207.645 97.430 ;
        RECT 208.235 97.340 208.420 97.430 ;
        RECT 203.580 96.380 203.870 97.050 ;
        RECT 204.050 96.560 204.515 96.870 ;
        RECT 204.695 96.560 205.220 96.870 ;
        RECT 203.580 96.180 204.810 96.380 ;
        RECT 203.650 95.630 204.320 96.000 ;
        RECT 204.500 95.810 204.810 96.180 ;
        RECT 204.990 95.920 205.220 96.560 ;
        RECT 205.400 96.540 205.700 96.870 ;
        RECT 205.400 95.630 205.690 96.360 ;
        RECT 205.880 96.140 206.050 97.330 ;
        RECT 207.750 97.230 208.080 97.260 ;
        RECT 206.280 97.170 208.080 97.230 ;
        RECT 208.670 97.170 208.925 97.790 ;
        RECT 209.215 97.550 209.500 98.010 ;
        RECT 209.670 97.720 209.940 98.180 ;
        RECT 209.215 97.330 210.170 97.550 ;
        RECT 206.220 97.060 208.925 97.170 ;
        RECT 206.220 97.025 206.420 97.060 ;
        RECT 206.220 96.450 206.390 97.025 ;
        RECT 207.750 97.000 208.925 97.060 ;
        RECT 206.620 96.585 207.030 96.890 ;
        RECT 207.200 96.620 207.530 96.830 ;
        RECT 206.220 96.330 206.490 96.450 ;
        RECT 206.220 96.285 207.065 96.330 ;
        RECT 206.310 96.160 207.065 96.285 ;
        RECT 207.320 96.220 207.530 96.620 ;
        RECT 207.775 96.620 208.250 96.830 ;
        RECT 208.440 96.620 208.930 96.820 ;
        RECT 207.775 96.220 207.995 96.620 ;
        RECT 209.100 96.600 209.790 97.160 ;
        RECT 209.960 96.430 210.170 97.330 ;
        RECT 205.880 96.130 206.110 96.140 ;
        RECT 205.880 95.800 206.140 96.130 ;
        RECT 206.895 96.010 207.065 96.160 ;
        RECT 206.310 95.630 206.640 95.990 ;
        RECT 206.895 95.800 208.195 96.010 ;
        RECT 208.470 95.630 208.925 96.395 ;
        RECT 209.215 96.260 210.170 96.430 ;
        RECT 210.340 97.160 210.740 98.010 ;
        RECT 210.930 97.550 211.210 98.010 ;
        RECT 211.730 97.720 212.055 98.180 ;
        RECT 210.930 97.330 212.055 97.550 ;
        RECT 210.340 96.600 211.435 97.160 ;
        RECT 211.605 96.870 212.055 97.330 ;
        RECT 212.225 97.040 212.610 98.010 ;
        RECT 212.780 97.745 218.125 98.180 ;
        RECT 209.215 95.800 209.500 96.260 ;
        RECT 209.670 95.630 209.940 96.090 ;
        RECT 210.340 95.800 210.740 96.600 ;
        RECT 211.605 96.540 212.160 96.870 ;
        RECT 211.605 96.430 212.055 96.540 ;
        RECT 210.930 96.260 212.055 96.430 ;
        RECT 212.330 96.370 212.610 97.040 ;
        RECT 210.930 95.800 211.210 96.260 ;
        RECT 211.730 95.630 212.055 96.090 ;
        RECT 212.225 95.800 212.610 96.370 ;
        RECT 214.365 96.175 214.705 97.005 ;
        RECT 216.185 96.495 216.535 97.745 ;
        RECT 218.300 97.090 221.810 98.180 ;
        RECT 221.980 97.090 223.190 98.180 ;
        RECT 218.300 96.400 219.950 96.920 ;
        RECT 220.120 96.570 221.810 97.090 ;
        RECT 212.780 95.630 218.125 96.175 ;
        RECT 218.300 95.630 221.810 96.400 ;
        RECT 221.980 96.380 222.500 96.920 ;
        RECT 222.670 96.550 223.190 97.090 ;
        RECT 223.365 97.790 223.700 98.010 ;
        RECT 224.705 97.800 225.060 98.180 ;
        RECT 223.365 97.170 223.620 97.790 ;
        RECT 223.870 97.630 224.100 97.670 ;
        RECT 225.230 97.630 225.480 98.010 ;
        RECT 223.870 97.430 225.480 97.630 ;
        RECT 223.870 97.340 224.055 97.430 ;
        RECT 224.645 97.420 225.480 97.430 ;
        RECT 225.730 97.400 225.980 98.180 ;
        RECT 226.150 97.330 226.410 98.010 ;
        RECT 224.210 97.230 224.540 97.260 ;
        RECT 224.210 97.170 226.010 97.230 ;
        RECT 223.365 97.060 226.070 97.170 ;
        RECT 223.365 97.000 224.540 97.060 ;
        RECT 225.870 97.025 226.070 97.060 ;
        RECT 223.360 96.620 223.850 96.820 ;
        RECT 224.040 96.620 224.515 96.830 ;
        RECT 221.980 95.630 223.190 96.380 ;
        RECT 223.365 95.630 223.820 96.395 ;
        RECT 224.295 96.220 224.515 96.620 ;
        RECT 224.760 96.620 225.090 96.830 ;
        RECT 224.760 96.220 224.970 96.620 ;
        RECT 225.260 96.585 225.670 96.890 ;
        RECT 225.900 96.450 226.070 97.025 ;
        RECT 225.800 96.330 226.070 96.450 ;
        RECT 225.225 96.285 226.070 96.330 ;
        RECT 225.225 96.160 225.980 96.285 ;
        RECT 225.225 96.010 225.395 96.160 ;
        RECT 226.240 96.130 226.410 97.330 ;
        RECT 226.580 97.015 226.870 98.180 ;
        RECT 227.590 97.170 227.760 98.010 ;
        RECT 227.930 97.840 229.100 98.010 ;
        RECT 227.930 97.340 228.260 97.840 ;
        RECT 228.770 97.800 229.100 97.840 ;
        RECT 229.290 97.760 229.645 98.180 ;
        RECT 228.430 97.580 228.660 97.670 ;
        RECT 229.815 97.580 230.065 98.010 ;
        RECT 228.430 97.340 230.065 97.580 ;
        RECT 230.235 97.420 230.565 98.180 ;
        RECT 230.735 97.340 230.990 98.010 ;
        RECT 231.180 97.745 236.525 98.180 ;
        RECT 227.590 97.000 230.650 97.170 ;
        RECT 227.505 96.620 227.855 96.830 ;
        RECT 228.025 96.620 228.470 96.820 ;
        RECT 228.640 96.620 229.115 96.820 ;
        RECT 224.095 95.800 225.395 96.010 ;
        RECT 225.650 95.630 225.980 95.990 ;
        RECT 226.150 95.800 226.410 96.130 ;
        RECT 226.580 95.630 226.870 96.355 ;
        RECT 227.590 96.280 228.655 96.450 ;
        RECT 227.590 95.800 227.760 96.280 ;
        RECT 227.930 95.630 228.260 96.110 ;
        RECT 228.485 96.050 228.655 96.280 ;
        RECT 228.835 96.220 229.115 96.620 ;
        RECT 229.385 96.620 229.715 96.820 ;
        RECT 229.885 96.650 230.260 96.820 ;
        RECT 229.885 96.620 230.250 96.650 ;
        RECT 229.385 96.220 229.670 96.620 ;
        RECT 230.480 96.450 230.650 97.000 ;
        RECT 229.850 96.280 230.650 96.450 ;
        RECT 229.850 96.050 230.020 96.280 ;
        RECT 230.820 96.210 230.990 97.340 ;
        RECT 230.805 96.140 230.990 96.210 ;
        RECT 232.765 96.175 233.105 97.005 ;
        RECT 234.585 96.495 234.935 97.745 ;
        RECT 236.700 97.090 240.210 98.180 ;
        RECT 236.700 96.400 238.350 96.920 ;
        RECT 238.520 96.570 240.210 97.090 ;
        RECT 240.840 97.330 241.100 98.010 ;
        RECT 241.270 97.400 241.520 98.180 ;
        RECT 241.770 97.630 242.020 98.010 ;
        RECT 242.190 97.800 242.545 98.180 ;
        RECT 243.550 97.790 243.885 98.010 ;
        RECT 243.150 97.630 243.380 97.670 ;
        RECT 241.770 97.430 243.380 97.630 ;
        RECT 241.770 97.420 242.605 97.430 ;
        RECT 243.195 97.340 243.380 97.430 ;
        RECT 230.780 96.130 230.990 96.140 ;
        RECT 228.485 95.800 230.020 96.050 ;
        RECT 230.190 95.630 230.520 96.110 ;
        RECT 230.735 95.800 230.990 96.130 ;
        RECT 231.180 95.630 236.525 96.175 ;
        RECT 236.700 95.630 240.210 96.400 ;
        RECT 240.840 96.130 241.010 97.330 ;
        RECT 242.710 97.230 243.040 97.260 ;
        RECT 241.240 97.170 243.040 97.230 ;
        RECT 243.630 97.170 243.885 97.790 ;
        RECT 241.180 97.060 243.885 97.170 ;
        RECT 241.180 97.025 241.380 97.060 ;
        RECT 241.180 96.450 241.350 97.025 ;
        RECT 242.710 97.000 243.885 97.060 ;
        RECT 244.065 97.790 244.400 98.010 ;
        RECT 245.405 97.800 245.760 98.180 ;
        RECT 244.065 97.170 244.320 97.790 ;
        RECT 244.570 97.630 244.800 97.670 ;
        RECT 245.930 97.630 246.180 98.010 ;
        RECT 244.570 97.430 246.180 97.630 ;
        RECT 244.570 97.340 244.755 97.430 ;
        RECT 245.345 97.420 246.180 97.430 ;
        RECT 246.430 97.400 246.680 98.180 ;
        RECT 246.850 97.330 247.110 98.010 ;
        RECT 244.910 97.230 245.240 97.260 ;
        RECT 244.910 97.170 246.710 97.230 ;
        RECT 244.065 97.060 246.770 97.170 ;
        RECT 244.065 97.000 245.240 97.060 ;
        RECT 246.570 97.025 246.770 97.060 ;
        RECT 241.580 96.585 241.990 96.890 ;
        RECT 242.160 96.620 242.490 96.830 ;
        RECT 241.180 96.330 241.450 96.450 ;
        RECT 241.180 96.285 242.025 96.330 ;
        RECT 241.270 96.160 242.025 96.285 ;
        RECT 242.280 96.220 242.490 96.620 ;
        RECT 242.735 96.620 243.210 96.830 ;
        RECT 243.400 96.620 243.890 96.820 ;
        RECT 244.060 96.620 244.550 96.820 ;
        RECT 244.740 96.620 245.215 96.830 ;
        RECT 242.735 96.220 242.955 96.620 ;
        RECT 240.840 95.800 241.100 96.130 ;
        RECT 241.855 96.010 242.025 96.160 ;
        RECT 241.270 95.630 241.600 95.990 ;
        RECT 241.855 95.800 243.155 96.010 ;
        RECT 243.430 95.630 243.885 96.395 ;
        RECT 244.065 95.630 244.520 96.395 ;
        RECT 244.995 96.220 245.215 96.620 ;
        RECT 245.460 96.620 245.790 96.830 ;
        RECT 245.460 96.220 245.670 96.620 ;
        RECT 245.960 96.585 246.370 96.890 ;
        RECT 246.600 96.450 246.770 97.025 ;
        RECT 246.500 96.330 246.770 96.450 ;
        RECT 245.925 96.285 246.770 96.330 ;
        RECT 245.925 96.160 246.680 96.285 ;
        RECT 245.925 96.010 246.095 96.160 ;
        RECT 246.940 96.140 247.110 97.330 ;
        RECT 246.880 96.130 247.110 96.140 ;
        RECT 244.795 95.800 246.095 96.010 ;
        RECT 246.350 95.630 246.680 95.990 ;
        RECT 246.850 95.800 247.110 96.130 ;
        RECT 248.220 97.340 248.475 98.010 ;
        RECT 248.645 97.420 248.975 98.180 ;
        RECT 249.145 97.580 249.395 98.010 ;
        RECT 249.565 97.760 249.920 98.180 ;
        RECT 250.110 97.840 251.280 98.010 ;
        RECT 250.110 97.800 250.440 97.840 ;
        RECT 250.550 97.580 250.780 97.670 ;
        RECT 249.145 97.340 250.780 97.580 ;
        RECT 250.950 97.340 251.280 97.840 ;
        RECT 248.220 97.330 248.430 97.340 ;
        RECT 248.220 96.210 248.390 97.330 ;
        RECT 251.450 97.170 251.620 98.010 ;
        RECT 248.560 97.000 251.620 97.170 ;
        RECT 252.340 97.015 252.630 98.180 ;
        RECT 252.800 97.330 253.060 98.010 ;
        RECT 253.230 97.400 253.480 98.180 ;
        RECT 253.730 97.630 253.980 98.010 ;
        RECT 254.150 97.800 254.505 98.180 ;
        RECT 255.510 97.790 255.845 98.010 ;
        RECT 255.110 97.630 255.340 97.670 ;
        RECT 253.730 97.430 255.340 97.630 ;
        RECT 253.730 97.420 254.565 97.430 ;
        RECT 255.155 97.340 255.340 97.430 ;
        RECT 248.560 96.450 248.730 97.000 ;
        RECT 248.960 96.620 249.325 96.820 ;
        RECT 249.495 96.620 249.825 96.820 ;
        RECT 248.560 96.280 249.360 96.450 ;
        RECT 248.220 96.130 248.405 96.210 ;
        RECT 248.220 95.800 248.475 96.130 ;
        RECT 248.690 95.630 249.020 96.110 ;
        RECT 249.190 96.050 249.360 96.280 ;
        RECT 249.540 96.220 249.825 96.620 ;
        RECT 250.095 96.620 250.570 96.820 ;
        RECT 250.740 96.620 251.185 96.820 ;
        RECT 251.355 96.620 251.705 96.830 ;
        RECT 250.095 96.220 250.375 96.620 ;
        RECT 250.555 96.280 251.620 96.450 ;
        RECT 250.555 96.050 250.725 96.280 ;
        RECT 249.190 95.800 250.725 96.050 ;
        RECT 250.950 95.630 251.280 96.110 ;
        RECT 251.450 95.800 251.620 96.280 ;
        RECT 252.340 95.630 252.630 96.355 ;
        RECT 252.800 96.130 252.970 97.330 ;
        RECT 254.670 97.230 255.000 97.260 ;
        RECT 253.200 97.170 255.000 97.230 ;
        RECT 255.590 97.170 255.845 97.790 ;
        RECT 253.140 97.060 255.845 97.170 ;
        RECT 256.030 97.115 256.340 98.180 ;
        RECT 256.510 97.510 256.745 98.010 ;
        RECT 256.915 97.720 257.245 98.180 ;
        RECT 257.440 97.840 258.550 98.010 ;
        RECT 257.440 97.680 257.630 97.840 ;
        RECT 257.860 97.510 258.160 97.670 ;
        RECT 256.510 97.330 258.160 97.510 ;
        RECT 258.330 97.330 258.550 97.840 ;
        RECT 258.720 97.330 259.050 98.180 ;
        RECT 259.240 97.745 264.585 98.180 ;
        RECT 253.140 97.025 253.340 97.060 ;
        RECT 253.140 96.450 253.310 97.025 ;
        RECT 254.670 97.000 255.845 97.060 ;
        RECT 253.540 96.585 253.950 96.890 ;
        RECT 254.120 96.620 254.450 96.830 ;
        RECT 253.140 96.330 253.410 96.450 ;
        RECT 253.140 96.285 253.985 96.330 ;
        RECT 253.230 96.160 253.985 96.285 ;
        RECT 254.240 96.220 254.450 96.620 ;
        RECT 254.695 96.620 255.170 96.830 ;
        RECT 255.360 96.620 255.850 96.820 ;
        RECT 254.695 96.220 254.915 96.620 ;
        RECT 252.800 95.800 253.060 96.130 ;
        RECT 253.815 96.010 253.985 96.160 ;
        RECT 253.230 95.630 253.560 95.990 ;
        RECT 253.815 95.800 255.115 96.010 ;
        RECT 255.390 95.630 255.845 96.395 ;
        RECT 256.025 96.310 256.340 96.945 ;
        RECT 256.510 96.140 256.720 97.330 ;
        RECT 257.060 96.990 259.035 97.160 ;
        RECT 257.060 96.620 257.555 96.990 ;
        RECT 257.735 96.620 258.535 96.820 ;
        RECT 258.705 96.600 259.035 96.990 ;
        RECT 256.890 96.260 259.050 96.430 ;
        RECT 256.030 95.970 256.340 96.140 ;
        RECT 256.890 95.970 257.220 96.260 ;
        RECT 256.030 95.800 257.220 95.970 ;
        RECT 257.460 95.630 257.630 96.090 ;
        RECT 257.860 95.800 258.190 96.260 ;
        RECT 258.370 95.630 258.540 96.090 ;
        RECT 258.720 95.800 259.050 96.260 ;
        RECT 260.825 96.175 261.165 97.005 ;
        RECT 262.645 96.495 262.995 97.745 ;
        RECT 264.760 97.090 268.270 98.180 ;
        RECT 264.760 96.400 266.410 96.920 ;
        RECT 266.580 96.570 268.270 97.090 ;
        RECT 269.365 97.030 269.625 98.180 ;
        RECT 269.800 97.105 270.055 98.010 ;
        RECT 270.225 97.420 270.555 98.180 ;
        RECT 270.770 97.250 270.940 98.010 ;
        RECT 259.240 95.630 264.585 96.175 ;
        RECT 264.760 95.630 268.270 96.400 ;
        RECT 269.365 95.630 269.625 96.470 ;
        RECT 269.800 96.375 269.970 97.105 ;
        RECT 270.225 97.080 270.940 97.250 ;
        RECT 270.225 96.870 270.395 97.080 ;
        RECT 271.205 97.030 271.465 98.180 ;
        RECT 271.640 97.105 271.895 98.010 ;
        RECT 272.065 97.420 272.395 98.180 ;
        RECT 272.610 97.250 272.780 98.010 ;
        RECT 270.140 96.540 270.395 96.870 ;
        RECT 269.800 95.800 270.055 96.375 ;
        RECT 270.225 96.350 270.395 96.540 ;
        RECT 270.675 96.530 271.030 96.900 ;
        RECT 270.225 96.180 270.940 96.350 ;
        RECT 270.225 95.630 270.555 96.010 ;
        RECT 270.770 95.800 270.940 96.180 ;
        RECT 271.205 95.630 271.465 96.470 ;
        RECT 271.640 96.375 271.810 97.105 ;
        RECT 272.065 97.080 272.780 97.250 ;
        RECT 272.065 96.870 272.235 97.080 ;
        RECT 273.965 97.040 274.300 98.010 ;
        RECT 274.470 97.040 274.640 98.180 ;
        RECT 274.810 97.840 276.840 98.010 ;
        RECT 271.980 96.540 272.235 96.870 ;
        RECT 271.640 95.800 271.895 96.375 ;
        RECT 272.065 96.350 272.235 96.540 ;
        RECT 272.515 96.530 272.870 96.900 ;
        RECT 273.965 96.370 274.135 97.040 ;
        RECT 274.810 96.870 274.980 97.840 ;
        RECT 274.305 96.540 274.560 96.870 ;
        RECT 274.785 96.540 274.980 96.870 ;
        RECT 275.150 97.500 276.275 97.670 ;
        RECT 274.390 96.370 274.560 96.540 ;
        RECT 275.150 96.370 275.320 97.500 ;
        RECT 272.065 96.180 272.780 96.350 ;
        RECT 272.065 95.630 272.395 96.010 ;
        RECT 272.610 95.800 272.780 96.180 ;
        RECT 273.965 95.800 274.220 96.370 ;
        RECT 274.390 96.200 275.320 96.370 ;
        RECT 275.490 97.160 276.500 97.330 ;
        RECT 275.490 96.360 275.660 97.160 ;
        RECT 275.145 96.165 275.320 96.200 ;
        RECT 274.390 95.630 274.720 96.030 ;
        RECT 275.145 95.800 275.675 96.165 ;
        RECT 275.865 96.140 276.140 96.960 ;
        RECT 275.860 95.970 276.140 96.140 ;
        RECT 275.865 95.800 276.140 95.970 ;
        RECT 276.310 95.800 276.500 97.160 ;
        RECT 276.670 97.175 276.840 97.840 ;
        RECT 277.010 97.420 277.180 98.180 ;
        RECT 277.415 97.420 277.930 97.830 ;
        RECT 276.670 96.985 277.420 97.175 ;
        RECT 277.590 96.610 277.930 97.420 ;
        RECT 278.100 97.015 278.390 98.180 ;
        RECT 278.560 97.420 279.075 97.830 ;
        RECT 279.310 97.420 279.480 98.180 ;
        RECT 279.650 97.840 281.680 98.010 ;
        RECT 276.700 96.440 277.930 96.610 ;
        RECT 278.560 96.610 278.900 97.420 ;
        RECT 279.650 97.175 279.820 97.840 ;
        RECT 280.215 97.500 281.340 97.670 ;
        RECT 279.070 96.985 279.820 97.175 ;
        RECT 279.990 97.160 281.000 97.330 ;
        RECT 278.560 96.440 279.790 96.610 ;
        RECT 276.680 95.630 277.190 96.165 ;
        RECT 277.410 95.835 277.655 96.440 ;
        RECT 278.100 95.630 278.390 96.355 ;
        RECT 278.835 95.835 279.080 96.440 ;
        RECT 279.300 95.630 279.810 96.165 ;
        RECT 279.990 95.800 280.180 97.160 ;
        RECT 280.350 96.820 280.625 96.960 ;
        RECT 280.350 96.650 280.630 96.820 ;
        RECT 280.350 95.800 280.625 96.650 ;
        RECT 280.830 96.360 281.000 97.160 ;
        RECT 281.170 96.370 281.340 97.500 ;
        RECT 281.510 96.870 281.680 97.840 ;
        RECT 281.850 97.040 282.020 98.180 ;
        RECT 282.190 97.040 282.525 98.010 ;
        RECT 282.710 97.460 283.040 98.180 ;
        RECT 281.510 96.540 281.705 96.870 ;
        RECT 281.930 96.540 282.185 96.870 ;
        RECT 281.930 96.370 282.100 96.540 ;
        RECT 282.355 96.370 282.525 97.040 ;
        RECT 282.700 96.820 282.930 97.160 ;
        RECT 283.220 96.820 283.435 97.935 ;
        RECT 283.630 97.235 283.960 98.010 ;
        RECT 284.130 97.405 284.840 98.180 ;
        RECT 283.630 97.020 284.780 97.235 ;
        RECT 282.700 96.620 283.030 96.820 ;
        RECT 283.220 96.640 283.670 96.820 ;
        RECT 283.340 96.620 283.670 96.640 ;
        RECT 283.840 96.620 284.310 96.850 ;
        RECT 284.495 96.450 284.780 97.020 ;
        RECT 285.010 96.575 285.290 98.010 ;
        RECT 285.550 97.250 285.720 98.010 ;
        RECT 285.935 97.420 286.265 98.180 ;
        RECT 285.550 97.080 286.265 97.250 ;
        RECT 286.435 97.105 286.690 98.010 ;
        RECT 281.170 96.200 282.100 96.370 ;
        RECT 281.170 96.165 281.345 96.200 ;
        RECT 280.815 95.800 281.345 96.165 ;
        RECT 281.770 95.630 282.100 96.030 ;
        RECT 282.270 95.800 282.525 96.370 ;
        RECT 282.700 96.260 283.880 96.450 ;
        RECT 282.700 95.800 283.040 96.260 ;
        RECT 283.550 96.180 283.880 96.260 ;
        RECT 284.070 96.260 284.780 96.450 ;
        RECT 284.070 96.120 284.370 96.260 ;
        RECT 284.055 96.110 284.370 96.120 ;
        RECT 284.045 96.100 284.370 96.110 ;
        RECT 284.035 96.095 284.370 96.100 ;
        RECT 283.210 95.630 283.380 96.090 ;
        RECT 284.030 96.085 284.370 96.095 ;
        RECT 284.025 96.080 284.370 96.085 ;
        RECT 284.020 96.070 284.370 96.080 ;
        RECT 284.015 96.065 284.370 96.070 ;
        RECT 284.010 95.800 284.370 96.065 ;
        RECT 284.610 95.630 284.780 96.090 ;
        RECT 284.950 95.800 285.290 96.575 ;
        RECT 285.460 96.530 285.815 96.900 ;
        RECT 286.095 96.870 286.265 97.080 ;
        RECT 286.095 96.540 286.350 96.870 ;
        RECT 286.095 96.350 286.265 96.540 ;
        RECT 286.520 96.375 286.690 97.105 ;
        RECT 286.865 97.030 287.125 98.180 ;
        RECT 287.300 97.090 288.510 98.180 ;
        RECT 285.550 96.180 286.265 96.350 ;
        RECT 285.550 95.800 285.720 96.180 ;
        RECT 285.935 95.630 286.265 96.010 ;
        RECT 286.435 95.800 286.690 96.375 ;
        RECT 286.865 95.630 287.125 96.470 ;
        RECT 287.300 96.380 287.820 96.920 ;
        RECT 287.990 96.550 288.510 97.090 ;
        RECT 288.770 97.250 288.940 98.010 ;
        RECT 289.155 97.420 289.485 98.180 ;
        RECT 288.770 97.080 289.485 97.250 ;
        RECT 289.655 97.105 289.910 98.010 ;
        RECT 288.680 96.530 289.035 96.900 ;
        RECT 289.315 96.870 289.485 97.080 ;
        RECT 289.315 96.540 289.570 96.870 ;
        RECT 287.300 95.630 288.510 96.380 ;
        RECT 289.315 96.350 289.485 96.540 ;
        RECT 289.740 96.375 289.910 97.105 ;
        RECT 290.085 97.030 290.345 98.180 ;
        RECT 290.525 97.030 290.785 98.180 ;
        RECT 290.960 97.105 291.215 98.010 ;
        RECT 291.385 97.420 291.715 98.180 ;
        RECT 291.930 97.250 292.100 98.010 ;
        RECT 288.770 96.180 289.485 96.350 ;
        RECT 288.770 95.800 288.940 96.180 ;
        RECT 289.155 95.630 289.485 96.010 ;
        RECT 289.655 95.800 289.910 96.375 ;
        RECT 290.085 95.630 290.345 96.470 ;
        RECT 290.525 95.630 290.785 96.470 ;
        RECT 290.960 96.375 291.130 97.105 ;
        RECT 291.385 97.080 292.100 97.250 ;
        RECT 292.360 97.090 294.030 98.180 ;
        RECT 294.665 97.510 294.920 98.010 ;
        RECT 295.090 97.680 295.420 98.180 ;
        RECT 294.665 97.340 295.415 97.510 ;
        RECT 291.385 96.870 291.555 97.080 ;
        RECT 291.300 96.540 291.555 96.870 ;
        RECT 290.960 95.800 291.215 96.375 ;
        RECT 291.385 96.350 291.555 96.540 ;
        RECT 291.835 96.530 292.190 96.900 ;
        RECT 292.360 96.400 293.110 96.920 ;
        RECT 293.280 96.570 294.030 97.090 ;
        RECT 294.665 96.520 295.015 97.170 ;
        RECT 291.385 96.180 292.100 96.350 ;
        RECT 291.385 95.630 291.715 96.010 ;
        RECT 291.930 95.800 292.100 96.180 ;
        RECT 292.360 95.630 294.030 96.400 ;
        RECT 295.185 96.350 295.415 97.340 ;
        RECT 294.665 96.180 295.415 96.350 ;
        RECT 294.665 95.890 294.920 96.180 ;
        RECT 295.090 95.630 295.420 96.010 ;
        RECT 295.590 95.890 295.760 98.010 ;
        RECT 295.930 97.210 296.255 97.995 ;
        RECT 296.425 97.720 296.675 98.180 ;
        RECT 296.845 97.680 297.095 98.010 ;
        RECT 297.310 97.680 297.990 98.010 ;
        RECT 296.845 97.550 297.015 97.680 ;
        RECT 296.620 97.380 297.015 97.550 ;
        RECT 295.990 96.160 296.450 97.210 ;
        RECT 296.620 96.020 296.790 97.380 ;
        RECT 297.185 97.120 297.650 97.510 ;
        RECT 296.960 96.310 297.310 96.930 ;
        RECT 297.480 96.530 297.650 97.120 ;
        RECT 297.820 96.900 297.990 97.680 ;
        RECT 298.160 97.580 298.330 97.920 ;
        RECT 298.565 97.750 298.895 98.180 ;
        RECT 299.065 97.580 299.235 97.920 ;
        RECT 299.530 97.720 299.900 98.180 ;
        RECT 298.160 97.410 299.235 97.580 ;
        RECT 300.070 97.550 300.240 98.010 ;
        RECT 300.475 97.670 301.345 98.010 ;
        RECT 301.515 97.720 301.765 98.180 ;
        RECT 299.680 97.380 300.240 97.550 ;
        RECT 299.680 97.240 299.850 97.380 ;
        RECT 298.350 97.070 299.850 97.240 ;
        RECT 300.545 97.210 301.005 97.500 ;
        RECT 297.820 96.730 299.510 96.900 ;
        RECT 297.480 96.310 297.835 96.530 ;
        RECT 298.005 96.020 298.175 96.730 ;
        RECT 298.380 96.310 299.170 96.560 ;
        RECT 299.340 96.550 299.510 96.730 ;
        RECT 299.680 96.380 299.850 97.070 ;
        RECT 296.120 95.630 296.450 95.990 ;
        RECT 296.620 95.850 297.115 96.020 ;
        RECT 297.320 95.850 298.175 96.020 ;
        RECT 299.050 95.630 299.380 96.090 ;
        RECT 299.590 95.990 299.850 96.380 ;
        RECT 300.040 97.200 301.005 97.210 ;
        RECT 301.175 97.290 301.345 97.670 ;
        RECT 301.935 97.630 302.105 97.920 ;
        RECT 302.285 97.800 302.615 98.180 ;
        RECT 301.935 97.460 302.735 97.630 ;
        RECT 300.040 97.040 300.715 97.200 ;
        RECT 301.175 97.120 302.395 97.290 ;
        RECT 300.040 96.250 300.250 97.040 ;
        RECT 301.175 97.030 301.345 97.120 ;
        RECT 300.420 96.250 300.770 96.870 ;
        RECT 300.940 96.860 301.345 97.030 ;
        RECT 300.940 96.080 301.110 96.860 ;
        RECT 301.280 96.410 301.500 96.690 ;
        RECT 301.680 96.580 302.220 96.950 ;
        RECT 302.565 96.870 302.735 97.460 ;
        RECT 302.955 97.040 303.260 98.180 ;
        RECT 303.430 96.990 303.685 97.870 ;
        RECT 303.860 97.015 304.150 98.180 ;
        RECT 304.325 97.040 304.660 98.010 ;
        RECT 304.830 97.040 305.000 98.180 ;
        RECT 305.170 97.840 307.200 98.010 ;
        RECT 302.565 96.840 303.305 96.870 ;
        RECT 301.280 96.240 301.810 96.410 ;
        RECT 299.590 95.820 299.940 95.990 ;
        RECT 300.160 95.800 301.110 96.080 ;
        RECT 301.280 95.630 301.470 96.070 ;
        RECT 301.640 96.010 301.810 96.240 ;
        RECT 301.980 96.180 302.220 96.580 ;
        RECT 302.390 96.540 303.305 96.840 ;
        RECT 302.390 96.365 302.715 96.540 ;
        RECT 302.390 96.010 302.710 96.365 ;
        RECT 303.475 96.340 303.685 96.990 ;
        RECT 304.325 96.370 304.495 97.040 ;
        RECT 305.170 96.870 305.340 97.840 ;
        RECT 304.665 96.540 304.920 96.870 ;
        RECT 305.145 96.540 305.340 96.870 ;
        RECT 305.510 97.500 306.635 97.670 ;
        RECT 304.750 96.370 304.920 96.540 ;
        RECT 305.510 96.370 305.680 97.500 ;
        RECT 301.640 95.840 302.710 96.010 ;
        RECT 302.955 95.630 303.260 96.090 ;
        RECT 303.430 95.810 303.685 96.340 ;
        RECT 303.860 95.630 304.150 96.355 ;
        RECT 304.325 95.800 304.580 96.370 ;
        RECT 304.750 96.200 305.680 96.370 ;
        RECT 305.850 97.160 306.860 97.330 ;
        RECT 305.850 96.360 306.020 97.160 ;
        RECT 305.505 96.165 305.680 96.200 ;
        RECT 304.750 95.630 305.080 96.030 ;
        RECT 305.505 95.800 306.035 96.165 ;
        RECT 306.225 96.140 306.500 96.960 ;
        RECT 306.220 95.970 306.500 96.140 ;
        RECT 306.225 95.800 306.500 95.970 ;
        RECT 306.670 95.800 306.860 97.160 ;
        RECT 307.030 97.175 307.200 97.840 ;
        RECT 307.370 97.420 307.540 98.180 ;
        RECT 307.775 97.420 308.290 97.830 ;
        RECT 307.030 96.985 307.780 97.175 ;
        RECT 307.950 96.610 308.290 97.420 ;
        RECT 308.460 97.090 309.670 98.180 ;
        RECT 307.060 96.440 308.290 96.610 ;
        RECT 307.040 95.630 307.550 96.165 ;
        RECT 307.770 95.835 308.015 96.440 ;
        RECT 308.460 96.380 308.980 96.920 ;
        RECT 309.150 96.550 309.670 97.090 ;
        RECT 309.840 97.090 311.050 98.180 ;
        RECT 309.840 96.550 310.360 97.090 ;
        RECT 310.530 96.380 311.050 96.920 ;
        RECT 308.460 95.630 309.670 96.380 ;
        RECT 309.840 95.630 311.050 96.380 ;
        RECT 162.095 95.460 311.135 95.630 ;
        RECT 162.180 94.710 163.390 95.460 ;
        RECT 162.180 94.170 162.700 94.710 ;
        RECT 163.565 94.620 163.825 95.460 ;
        RECT 164.000 94.715 164.255 95.290 ;
        RECT 164.425 95.080 164.755 95.460 ;
        RECT 164.970 94.910 165.140 95.290 ;
        RECT 164.425 94.740 165.140 94.910 ;
        RECT 162.870 94.000 163.390 94.540 ;
        RECT 162.180 92.910 163.390 94.000 ;
        RECT 163.565 92.910 163.825 94.060 ;
        RECT 164.000 93.985 164.170 94.715 ;
        RECT 164.425 94.550 164.595 94.740 ;
        RECT 165.400 94.690 168.910 95.460 ;
        RECT 169.080 94.710 170.290 95.460 ;
        RECT 170.465 94.910 170.720 95.200 ;
        RECT 170.890 95.080 171.220 95.460 ;
        RECT 170.465 94.740 171.215 94.910 ;
        RECT 164.340 94.220 164.595 94.550 ;
        RECT 164.425 94.010 164.595 94.220 ;
        RECT 164.875 94.190 165.230 94.560 ;
        RECT 165.400 94.170 167.050 94.690 ;
        RECT 164.000 93.080 164.255 93.985 ;
        RECT 164.425 93.840 165.140 94.010 ;
        RECT 167.220 94.000 168.910 94.520 ;
        RECT 169.080 94.170 169.600 94.710 ;
        RECT 169.770 94.000 170.290 94.540 ;
        RECT 164.425 92.910 164.755 93.670 ;
        RECT 164.970 93.080 165.140 93.840 ;
        RECT 165.400 92.910 168.910 94.000 ;
        RECT 169.080 92.910 170.290 94.000 ;
        RECT 170.465 93.920 170.815 94.570 ;
        RECT 170.985 93.750 171.215 94.740 ;
        RECT 170.465 93.580 171.215 93.750 ;
        RECT 170.465 93.080 170.720 93.580 ;
        RECT 170.890 92.910 171.220 93.410 ;
        RECT 171.390 93.080 171.560 95.200 ;
        RECT 171.920 95.100 172.250 95.460 ;
        RECT 172.420 95.070 172.915 95.240 ;
        RECT 173.120 95.070 173.975 95.240 ;
        RECT 171.790 93.880 172.250 94.930 ;
        RECT 171.730 93.095 172.055 93.880 ;
        RECT 172.420 93.710 172.590 95.070 ;
        RECT 172.760 94.160 173.110 94.780 ;
        RECT 173.280 94.560 173.635 94.780 ;
        RECT 173.280 93.970 173.450 94.560 ;
        RECT 173.805 94.360 173.975 95.070 ;
        RECT 174.850 95.000 175.180 95.460 ;
        RECT 175.390 95.100 175.740 95.270 ;
        RECT 174.180 94.530 174.970 94.780 ;
        RECT 175.390 94.710 175.650 95.100 ;
        RECT 175.960 95.010 176.910 95.290 ;
        RECT 177.080 95.020 177.270 95.460 ;
        RECT 177.440 95.080 178.510 95.250 ;
        RECT 175.140 94.360 175.310 94.540 ;
        RECT 172.420 93.540 172.815 93.710 ;
        RECT 172.985 93.580 173.450 93.970 ;
        RECT 173.620 94.190 175.310 94.360 ;
        RECT 172.645 93.410 172.815 93.540 ;
        RECT 173.620 93.410 173.790 94.190 ;
        RECT 175.480 94.020 175.650 94.710 ;
        RECT 174.150 93.850 175.650 94.020 ;
        RECT 175.840 94.050 176.050 94.840 ;
        RECT 176.220 94.220 176.570 94.840 ;
        RECT 176.740 94.230 176.910 95.010 ;
        RECT 177.440 94.850 177.610 95.080 ;
        RECT 177.080 94.680 177.610 94.850 ;
        RECT 177.080 94.400 177.300 94.680 ;
        RECT 177.780 94.510 178.020 94.910 ;
        RECT 176.740 94.060 177.145 94.230 ;
        RECT 177.480 94.140 178.020 94.510 ;
        RECT 178.190 94.725 178.510 95.080 ;
        RECT 178.755 95.000 179.060 95.460 ;
        RECT 179.230 94.750 179.485 95.280 ;
        RECT 179.660 94.915 185.005 95.460 ;
        RECT 178.190 94.550 178.515 94.725 ;
        RECT 178.190 94.250 179.105 94.550 ;
        RECT 178.365 94.220 179.105 94.250 ;
        RECT 175.840 93.890 176.515 94.050 ;
        RECT 176.975 93.970 177.145 94.060 ;
        RECT 175.840 93.880 176.805 93.890 ;
        RECT 175.480 93.710 175.650 93.850 ;
        RECT 172.225 92.910 172.475 93.370 ;
        RECT 172.645 93.080 172.895 93.410 ;
        RECT 173.110 93.080 173.790 93.410 ;
        RECT 173.960 93.510 175.035 93.680 ;
        RECT 175.480 93.540 176.040 93.710 ;
        RECT 176.345 93.590 176.805 93.880 ;
        RECT 176.975 93.800 178.195 93.970 ;
        RECT 173.960 93.170 174.130 93.510 ;
        RECT 174.365 92.910 174.695 93.340 ;
        RECT 174.865 93.170 175.035 93.510 ;
        RECT 175.330 92.910 175.700 93.370 ;
        RECT 175.870 93.080 176.040 93.540 ;
        RECT 176.975 93.420 177.145 93.800 ;
        RECT 178.365 93.630 178.535 94.220 ;
        RECT 179.275 94.100 179.485 94.750 ;
        RECT 176.275 93.080 177.145 93.420 ;
        RECT 177.735 93.460 178.535 93.630 ;
        RECT 177.315 92.910 177.565 93.370 ;
        RECT 177.735 93.170 177.905 93.460 ;
        RECT 178.085 92.910 178.415 93.290 ;
        RECT 178.755 92.910 179.060 94.050 ;
        RECT 179.230 93.220 179.485 94.100 ;
        RECT 181.245 94.085 181.585 94.915 ;
        RECT 185.180 94.690 187.770 95.460 ;
        RECT 187.940 94.735 188.230 95.460 ;
        RECT 189.320 94.960 189.620 95.290 ;
        RECT 189.790 94.980 190.065 95.460 ;
        RECT 183.065 93.345 183.415 94.595 ;
        RECT 185.180 94.170 186.390 94.690 ;
        RECT 186.560 94.000 187.770 94.520 ;
        RECT 179.660 92.910 185.005 93.345 ;
        RECT 185.180 92.910 187.770 94.000 ;
        RECT 187.940 92.910 188.230 94.075 ;
        RECT 189.320 94.050 189.490 94.960 ;
        RECT 190.245 94.810 190.540 95.200 ;
        RECT 190.710 94.980 190.965 95.460 ;
        RECT 191.140 94.810 191.400 95.200 ;
        RECT 191.570 94.980 191.850 95.460 ;
        RECT 189.660 94.220 190.010 94.790 ;
        RECT 190.245 94.640 191.895 94.810 ;
        RECT 190.180 94.300 191.320 94.470 ;
        RECT 190.180 94.050 190.350 94.300 ;
        RECT 191.490 94.130 191.895 94.640 ;
        RECT 189.320 93.880 190.350 94.050 ;
        RECT 191.140 93.960 191.895 94.130 ;
        RECT 192.080 94.515 192.420 95.290 ;
        RECT 192.590 95.000 192.760 95.460 ;
        RECT 193.000 95.025 193.360 95.290 ;
        RECT 193.000 95.020 193.355 95.025 ;
        RECT 193.000 95.010 193.350 95.020 ;
        RECT 193.000 95.005 193.345 95.010 ;
        RECT 193.000 94.995 193.340 95.005 ;
        RECT 193.990 95.000 194.160 95.460 ;
        RECT 193.000 94.990 193.335 94.995 ;
        RECT 193.000 94.980 193.325 94.990 ;
        RECT 193.000 94.970 193.315 94.980 ;
        RECT 193.000 94.830 193.300 94.970 ;
        RECT 192.590 94.640 193.300 94.830 ;
        RECT 193.490 94.830 193.820 94.910 ;
        RECT 194.330 94.830 194.670 95.290 ;
        RECT 194.840 94.915 200.185 95.460 ;
        RECT 200.360 94.915 205.705 95.460 ;
        RECT 193.490 94.640 194.670 94.830 ;
        RECT 189.320 93.080 189.630 93.880 ;
        RECT 191.140 93.710 191.400 93.960 ;
        RECT 189.800 92.910 190.110 93.710 ;
        RECT 190.280 93.540 191.400 93.710 ;
        RECT 190.280 93.080 190.540 93.540 ;
        RECT 190.710 92.910 190.965 93.370 ;
        RECT 191.140 93.080 191.400 93.540 ;
        RECT 191.570 92.910 191.855 93.780 ;
        RECT 192.080 93.080 192.360 94.515 ;
        RECT 192.590 94.070 192.875 94.640 ;
        RECT 193.060 94.240 193.530 94.470 ;
        RECT 193.700 94.450 194.030 94.470 ;
        RECT 193.700 94.270 194.150 94.450 ;
        RECT 194.340 94.270 194.670 94.470 ;
        RECT 192.590 93.855 193.740 94.070 ;
        RECT 192.530 92.910 193.240 93.685 ;
        RECT 193.410 93.080 193.740 93.855 ;
        RECT 193.935 93.155 194.150 94.270 ;
        RECT 194.440 93.930 194.670 94.270 ;
        RECT 196.425 94.085 196.765 94.915 ;
        RECT 194.330 92.910 194.660 93.630 ;
        RECT 198.245 93.345 198.595 94.595 ;
        RECT 201.945 94.085 202.285 94.915 ;
        RECT 203.765 93.345 204.115 94.595 ;
        RECT 194.840 92.910 200.185 93.345 ;
        RECT 200.360 92.910 205.705 93.345 ;
        RECT 205.890 93.090 206.150 95.280 ;
        RECT 206.410 95.090 207.080 95.460 ;
        RECT 207.260 94.910 207.570 95.280 ;
        RECT 206.340 94.710 207.570 94.910 ;
        RECT 206.340 94.040 206.630 94.710 ;
        RECT 207.750 94.530 207.980 95.170 ;
        RECT 208.160 94.730 208.450 95.460 ;
        RECT 208.645 94.695 209.100 95.460 ;
        RECT 209.375 95.080 210.675 95.290 ;
        RECT 210.930 95.100 211.260 95.460 ;
        RECT 210.505 94.930 210.675 95.080 ;
        RECT 211.430 94.960 211.690 95.290 ;
        RECT 206.810 94.220 207.275 94.530 ;
        RECT 207.455 94.220 207.980 94.530 ;
        RECT 208.160 94.220 208.460 94.550 ;
        RECT 209.575 94.470 209.795 94.870 ;
        RECT 208.640 94.270 209.130 94.470 ;
        RECT 209.320 94.260 209.795 94.470 ;
        RECT 210.040 94.470 210.250 94.870 ;
        RECT 210.505 94.805 211.260 94.930 ;
        RECT 210.505 94.760 211.350 94.805 ;
        RECT 211.080 94.640 211.350 94.760 ;
        RECT 210.040 94.260 210.370 94.470 ;
        RECT 210.540 94.200 210.950 94.505 ;
        RECT 206.340 93.820 207.110 94.040 ;
        RECT 206.320 92.910 206.660 93.640 ;
        RECT 206.840 93.090 207.110 93.820 ;
        RECT 207.290 93.800 208.450 94.040 ;
        RECT 207.290 93.090 207.520 93.800 ;
        RECT 207.690 92.910 208.020 93.620 ;
        RECT 208.190 93.090 208.450 93.800 ;
        RECT 208.645 94.030 209.820 94.090 ;
        RECT 211.180 94.065 211.350 94.640 ;
        RECT 211.150 94.030 211.350 94.065 ;
        RECT 208.645 93.920 211.350 94.030 ;
        RECT 208.645 93.300 208.900 93.920 ;
        RECT 209.490 93.860 211.290 93.920 ;
        RECT 209.490 93.830 209.820 93.860 ;
        RECT 211.520 93.760 211.690 94.960 ;
        RECT 211.860 94.690 213.530 95.460 ;
        RECT 213.700 94.735 213.990 95.460 ;
        RECT 214.160 94.915 219.505 95.460 ;
        RECT 219.680 94.915 225.025 95.460 ;
        RECT 226.140 94.960 226.395 95.290 ;
        RECT 226.610 94.980 226.940 95.460 ;
        RECT 227.110 95.040 228.645 95.290 ;
        RECT 226.140 94.950 226.350 94.960 ;
        RECT 211.860 94.170 212.610 94.690 ;
        RECT 212.780 94.000 213.530 94.520 ;
        RECT 215.745 94.085 216.085 94.915 ;
        RECT 209.150 93.660 209.335 93.750 ;
        RECT 209.925 93.660 210.760 93.670 ;
        RECT 209.150 93.460 210.760 93.660 ;
        RECT 209.150 93.420 209.380 93.460 ;
        RECT 208.645 93.080 208.980 93.300 ;
        RECT 209.985 92.910 210.340 93.290 ;
        RECT 210.510 93.080 210.760 93.460 ;
        RECT 211.010 92.910 211.260 93.690 ;
        RECT 211.430 93.080 211.690 93.760 ;
        RECT 211.860 92.910 213.530 94.000 ;
        RECT 213.700 92.910 213.990 94.075 ;
        RECT 217.565 93.345 217.915 94.595 ;
        RECT 221.265 94.085 221.605 94.915 ;
        RECT 226.140 94.880 226.325 94.950 ;
        RECT 223.085 93.345 223.435 94.595 ;
        RECT 226.140 93.750 226.310 94.880 ;
        RECT 227.110 94.810 227.280 95.040 ;
        RECT 226.480 94.640 227.280 94.810 ;
        RECT 226.480 94.090 226.650 94.640 ;
        RECT 227.460 94.470 227.745 94.870 ;
        RECT 226.880 94.440 227.245 94.470 ;
        RECT 226.870 94.270 227.245 94.440 ;
        RECT 227.415 94.270 227.745 94.470 ;
        RECT 228.015 94.470 228.295 94.870 ;
        RECT 228.475 94.810 228.645 95.040 ;
        RECT 228.870 94.980 229.200 95.460 ;
        RECT 229.370 94.810 229.540 95.290 ;
        RECT 229.800 94.915 235.145 95.460 ;
        RECT 228.475 94.640 229.540 94.810 ;
        RECT 228.015 94.270 228.490 94.470 ;
        RECT 228.660 94.270 229.105 94.470 ;
        RECT 229.275 94.260 229.625 94.470 ;
        RECT 226.480 93.920 229.540 94.090 ;
        RECT 231.385 94.085 231.725 94.915 ;
        RECT 235.320 94.690 238.830 95.460 ;
        RECT 239.460 94.735 239.750 95.460 ;
        RECT 239.920 94.710 241.130 95.460 ;
        RECT 241.320 94.960 241.575 95.290 ;
        RECT 241.790 94.980 242.120 95.460 ;
        RECT 242.290 95.040 243.825 95.290 ;
        RECT 241.320 94.880 241.505 94.960 ;
        RECT 214.160 92.910 219.505 93.345 ;
        RECT 219.680 92.910 225.025 93.345 ;
        RECT 226.140 93.080 226.395 93.750 ;
        RECT 226.565 92.910 226.895 93.670 ;
        RECT 227.065 93.510 228.700 93.750 ;
        RECT 227.065 93.080 227.315 93.510 ;
        RECT 228.470 93.420 228.700 93.510 ;
        RECT 227.485 92.910 227.840 93.330 ;
        RECT 228.030 93.250 228.360 93.290 ;
        RECT 228.870 93.250 229.200 93.750 ;
        RECT 228.030 93.080 229.200 93.250 ;
        RECT 229.370 93.080 229.540 93.920 ;
        RECT 233.205 93.345 233.555 94.595 ;
        RECT 235.320 94.170 236.970 94.690 ;
        RECT 237.140 94.000 238.830 94.520 ;
        RECT 239.920 94.170 240.440 94.710 ;
        RECT 229.800 92.910 235.145 93.345 ;
        RECT 235.320 92.910 238.830 94.000 ;
        RECT 239.460 92.910 239.750 94.075 ;
        RECT 240.610 94.000 241.130 94.540 ;
        RECT 239.920 92.910 241.130 94.000 ;
        RECT 241.320 93.760 241.490 94.880 ;
        RECT 242.290 94.810 242.460 95.040 ;
        RECT 241.660 94.640 242.460 94.810 ;
        RECT 241.660 94.090 241.830 94.640 ;
        RECT 242.640 94.470 242.925 94.870 ;
        RECT 242.060 94.270 242.425 94.470 ;
        RECT 242.595 94.270 242.925 94.470 ;
        RECT 243.195 94.470 243.475 94.870 ;
        RECT 243.655 94.810 243.825 95.040 ;
        RECT 244.050 94.980 244.380 95.460 ;
        RECT 244.550 94.810 244.720 95.290 ;
        RECT 243.655 94.640 244.720 94.810 ;
        RECT 244.980 94.690 246.650 95.460 ;
        RECT 246.910 94.810 247.080 95.290 ;
        RECT 247.250 94.980 247.580 95.460 ;
        RECT 247.805 95.040 249.340 95.290 ;
        RECT 247.805 94.810 247.975 95.040 ;
        RECT 243.195 94.270 243.670 94.470 ;
        RECT 243.840 94.270 244.285 94.470 ;
        RECT 244.455 94.260 244.805 94.470 ;
        RECT 244.980 94.170 245.730 94.690 ;
        RECT 246.910 94.640 247.975 94.810 ;
        RECT 241.660 93.920 244.720 94.090 ;
        RECT 245.900 94.000 246.650 94.520 ;
        RECT 248.155 94.470 248.435 94.870 ;
        RECT 246.825 94.260 247.175 94.470 ;
        RECT 247.345 94.270 247.790 94.470 ;
        RECT 247.960 94.270 248.435 94.470 ;
        RECT 248.705 94.470 248.990 94.870 ;
        RECT 249.170 94.810 249.340 95.040 ;
        RECT 249.510 94.980 249.840 95.460 ;
        RECT 250.055 94.960 250.310 95.290 ;
        RECT 250.100 94.950 250.310 94.960 ;
        RECT 250.125 94.880 250.310 94.950 ;
        RECT 249.170 94.640 249.970 94.810 ;
        RECT 248.705 94.270 249.035 94.470 ;
        RECT 249.205 94.270 249.570 94.470 ;
        RECT 249.800 94.090 249.970 94.640 ;
        RECT 241.320 93.750 241.530 93.760 ;
        RECT 241.320 93.080 241.575 93.750 ;
        RECT 241.745 92.910 242.075 93.670 ;
        RECT 242.245 93.510 243.880 93.750 ;
        RECT 242.245 93.080 242.495 93.510 ;
        RECT 243.650 93.420 243.880 93.510 ;
        RECT 242.665 92.910 243.020 93.330 ;
        RECT 243.210 93.250 243.540 93.290 ;
        RECT 244.050 93.250 244.380 93.750 ;
        RECT 243.210 93.080 244.380 93.250 ;
        RECT 244.550 93.080 244.720 93.920 ;
        RECT 244.980 92.910 246.650 94.000 ;
        RECT 246.910 93.920 249.970 94.090 ;
        RECT 246.910 93.080 247.080 93.920 ;
        RECT 250.140 93.750 250.310 94.880 ;
        RECT 247.250 93.250 247.580 93.750 ;
        RECT 247.750 93.510 249.385 93.750 ;
        RECT 247.750 93.420 247.980 93.510 ;
        RECT 248.090 93.250 248.420 93.290 ;
        RECT 247.250 93.080 248.420 93.250 ;
        RECT 248.610 92.910 248.965 93.330 ;
        RECT 249.135 93.080 249.385 93.510 ;
        RECT 249.555 92.910 249.885 93.670 ;
        RECT 250.055 93.080 250.310 93.750 ;
        RECT 250.520 94.960 250.775 95.290 ;
        RECT 250.990 94.980 251.320 95.460 ;
        RECT 251.490 95.040 253.025 95.290 ;
        RECT 250.520 94.880 250.705 94.960 ;
        RECT 250.520 93.750 250.690 94.880 ;
        RECT 251.490 94.810 251.660 95.040 ;
        RECT 250.860 94.640 251.660 94.810 ;
        RECT 250.860 94.090 251.030 94.640 ;
        RECT 251.840 94.470 252.125 94.870 ;
        RECT 251.260 94.270 251.625 94.470 ;
        RECT 251.795 94.270 252.125 94.470 ;
        RECT 252.395 94.470 252.675 94.870 ;
        RECT 252.855 94.810 253.025 95.040 ;
        RECT 253.250 94.980 253.580 95.460 ;
        RECT 253.750 94.810 253.920 95.290 ;
        RECT 254.180 94.915 259.525 95.460 ;
        RECT 259.700 94.915 265.045 95.460 ;
        RECT 252.855 94.640 253.920 94.810 ;
        RECT 252.395 94.270 252.870 94.470 ;
        RECT 253.040 94.270 253.485 94.470 ;
        RECT 253.655 94.260 254.005 94.470 ;
        RECT 250.860 93.920 253.920 94.090 ;
        RECT 255.765 94.085 256.105 94.915 ;
        RECT 250.520 93.080 250.775 93.750 ;
        RECT 250.945 92.910 251.275 93.670 ;
        RECT 251.445 93.510 253.080 93.750 ;
        RECT 251.445 93.080 251.695 93.510 ;
        RECT 252.850 93.420 253.080 93.510 ;
        RECT 251.865 92.910 252.220 93.330 ;
        RECT 252.410 93.250 252.740 93.290 ;
        RECT 253.250 93.250 253.580 93.750 ;
        RECT 252.410 93.080 253.580 93.250 ;
        RECT 253.750 93.080 253.920 93.920 ;
        RECT 257.585 93.345 257.935 94.595 ;
        RECT 261.285 94.085 261.625 94.915 ;
        RECT 265.220 94.735 265.510 95.460 ;
        RECT 265.680 94.915 271.025 95.460 ;
        RECT 271.200 94.915 276.545 95.460 ;
        RECT 263.105 93.345 263.455 94.595 ;
        RECT 267.265 94.085 267.605 94.915 ;
        RECT 254.180 92.910 259.525 93.345 ;
        RECT 259.700 92.910 265.045 93.345 ;
        RECT 265.220 92.910 265.510 94.075 ;
        RECT 269.085 93.345 269.435 94.595 ;
        RECT 272.785 94.085 273.125 94.915 ;
        RECT 277.180 94.830 277.520 95.290 ;
        RECT 277.690 95.000 277.860 95.460 ;
        RECT 278.490 95.025 278.850 95.290 ;
        RECT 278.495 95.020 278.850 95.025 ;
        RECT 278.500 95.010 278.850 95.020 ;
        RECT 278.505 95.005 278.850 95.010 ;
        RECT 278.510 94.995 278.850 95.005 ;
        RECT 279.090 95.000 279.260 95.460 ;
        RECT 278.515 94.990 278.850 94.995 ;
        RECT 278.525 94.980 278.850 94.990 ;
        RECT 278.535 94.970 278.850 94.980 ;
        RECT 278.030 94.830 278.360 94.910 ;
        RECT 277.180 94.640 278.360 94.830 ;
        RECT 278.550 94.830 278.850 94.970 ;
        RECT 278.550 94.640 279.260 94.830 ;
        RECT 274.605 93.345 274.955 94.595 ;
        RECT 277.180 94.270 277.510 94.470 ;
        RECT 277.820 94.450 278.150 94.470 ;
        RECT 277.700 94.270 278.150 94.450 ;
        RECT 277.180 93.930 277.410 94.270 ;
        RECT 265.680 92.910 271.025 93.345 ;
        RECT 271.200 92.910 276.545 93.345 ;
        RECT 277.190 92.910 277.520 93.630 ;
        RECT 277.700 93.155 277.915 94.270 ;
        RECT 278.320 94.240 278.790 94.470 ;
        RECT 278.975 94.070 279.260 94.640 ;
        RECT 279.430 94.515 279.770 95.290 ;
        RECT 278.110 93.855 279.260 94.070 ;
        RECT 278.110 93.080 278.440 93.855 ;
        RECT 278.610 92.910 279.320 93.685 ;
        RECT 279.490 93.080 279.770 94.515 ;
        RECT 279.940 94.690 281.610 95.460 ;
        RECT 281.780 94.830 282.120 95.290 ;
        RECT 282.290 95.000 282.460 95.460 ;
        RECT 283.090 95.025 283.450 95.290 ;
        RECT 283.095 95.020 283.450 95.025 ;
        RECT 283.100 95.010 283.450 95.020 ;
        RECT 283.105 95.005 283.450 95.010 ;
        RECT 283.110 94.995 283.450 95.005 ;
        RECT 283.690 95.000 283.860 95.460 ;
        RECT 283.115 94.990 283.450 94.995 ;
        RECT 283.125 94.980 283.450 94.990 ;
        RECT 283.135 94.970 283.450 94.980 ;
        RECT 282.630 94.830 282.960 94.910 ;
        RECT 279.940 94.170 280.690 94.690 ;
        RECT 281.780 94.640 282.960 94.830 ;
        RECT 283.150 94.830 283.450 94.970 ;
        RECT 283.150 94.640 283.860 94.830 ;
        RECT 280.860 94.000 281.610 94.520 ;
        RECT 279.940 92.910 281.610 94.000 ;
        RECT 281.780 94.270 282.110 94.470 ;
        RECT 282.420 94.450 282.750 94.470 ;
        RECT 282.300 94.270 282.750 94.450 ;
        RECT 281.780 93.930 282.010 94.270 ;
        RECT 281.790 92.910 282.120 93.630 ;
        RECT 282.300 93.155 282.515 94.270 ;
        RECT 282.920 94.240 283.390 94.470 ;
        RECT 283.575 94.070 283.860 94.640 ;
        RECT 284.030 94.515 284.370 95.290 ;
        RECT 284.540 94.915 289.885 95.460 ;
        RECT 282.710 93.855 283.860 94.070 ;
        RECT 282.710 93.080 283.040 93.855 ;
        RECT 283.210 92.910 283.920 93.685 ;
        RECT 284.090 93.080 284.370 94.515 ;
        RECT 286.125 94.085 286.465 94.915 ;
        RECT 290.980 94.735 291.270 95.460 ;
        RECT 291.445 94.720 291.700 95.290 ;
        RECT 291.870 95.060 292.200 95.460 ;
        RECT 292.625 94.925 293.155 95.290 ;
        RECT 292.625 94.890 292.800 94.925 ;
        RECT 291.870 94.720 292.800 94.890 ;
        RECT 287.945 93.345 288.295 94.595 ;
        RECT 284.540 92.910 289.885 93.345 ;
        RECT 290.980 92.910 291.270 94.075 ;
        RECT 291.445 94.050 291.615 94.720 ;
        RECT 291.870 94.550 292.040 94.720 ;
        RECT 291.785 94.220 292.040 94.550 ;
        RECT 292.265 94.220 292.460 94.550 ;
        RECT 291.445 93.080 291.780 94.050 ;
        RECT 291.950 92.910 292.120 94.050 ;
        RECT 292.290 93.250 292.460 94.220 ;
        RECT 292.630 93.590 292.800 94.720 ;
        RECT 292.970 93.930 293.140 94.730 ;
        RECT 293.345 94.440 293.620 95.290 ;
        RECT 293.340 94.270 293.620 94.440 ;
        RECT 293.345 94.130 293.620 94.270 ;
        RECT 293.790 93.930 293.980 95.290 ;
        RECT 294.160 94.925 294.670 95.460 ;
        RECT 294.890 94.650 295.135 95.255 ;
        RECT 296.505 94.720 296.760 95.290 ;
        RECT 296.930 95.060 297.260 95.460 ;
        RECT 297.685 94.925 298.215 95.290 ;
        RECT 298.405 95.120 298.680 95.290 ;
        RECT 298.400 94.950 298.680 95.120 ;
        RECT 297.685 94.890 297.860 94.925 ;
        RECT 296.930 94.720 297.860 94.890 ;
        RECT 294.180 94.480 295.410 94.650 ;
        RECT 292.970 93.760 293.980 93.930 ;
        RECT 294.150 93.915 294.900 94.105 ;
        RECT 292.630 93.420 293.755 93.590 ;
        RECT 294.150 93.250 294.320 93.915 ;
        RECT 295.070 93.670 295.410 94.480 ;
        RECT 292.290 93.080 294.320 93.250 ;
        RECT 294.490 92.910 294.660 93.670 ;
        RECT 294.895 93.260 295.410 93.670 ;
        RECT 296.505 94.050 296.675 94.720 ;
        RECT 296.930 94.550 297.100 94.720 ;
        RECT 296.845 94.220 297.100 94.550 ;
        RECT 297.325 94.220 297.520 94.550 ;
        RECT 296.505 93.080 296.840 94.050 ;
        RECT 297.010 92.910 297.180 94.050 ;
        RECT 297.350 93.250 297.520 94.220 ;
        RECT 297.690 93.590 297.860 94.720 ;
        RECT 298.030 93.930 298.200 94.730 ;
        RECT 298.405 94.130 298.680 94.950 ;
        RECT 298.850 93.930 299.040 95.290 ;
        RECT 299.220 94.925 299.730 95.460 ;
        RECT 299.950 94.650 300.195 95.255 ;
        RECT 300.645 94.720 300.900 95.290 ;
        RECT 301.070 95.060 301.400 95.460 ;
        RECT 301.825 94.925 302.355 95.290 ;
        RECT 301.825 94.890 302.000 94.925 ;
        RECT 301.070 94.720 302.000 94.890 ;
        RECT 299.240 94.480 300.470 94.650 ;
        RECT 298.030 93.760 299.040 93.930 ;
        RECT 299.210 93.915 299.960 94.105 ;
        RECT 297.690 93.420 298.815 93.590 ;
        RECT 299.210 93.250 299.380 93.915 ;
        RECT 300.130 93.670 300.470 94.480 ;
        RECT 297.350 93.080 299.380 93.250 ;
        RECT 299.550 92.910 299.720 93.670 ;
        RECT 299.955 93.260 300.470 93.670 ;
        RECT 300.645 94.050 300.815 94.720 ;
        RECT 301.070 94.550 301.240 94.720 ;
        RECT 300.985 94.220 301.240 94.550 ;
        RECT 301.465 94.220 301.660 94.550 ;
        RECT 300.645 93.080 300.980 94.050 ;
        RECT 301.150 92.910 301.320 94.050 ;
        RECT 301.490 93.250 301.660 94.220 ;
        RECT 301.830 93.590 302.000 94.720 ;
        RECT 302.170 93.930 302.340 94.730 ;
        RECT 302.545 94.440 302.820 95.290 ;
        RECT 302.540 94.270 302.820 94.440 ;
        RECT 302.545 94.130 302.820 94.270 ;
        RECT 302.990 93.930 303.180 95.290 ;
        RECT 303.360 94.925 303.870 95.460 ;
        RECT 304.090 94.650 304.335 95.255 ;
        RECT 304.870 94.910 305.040 95.290 ;
        RECT 305.255 95.080 305.585 95.460 ;
        RECT 304.870 94.740 305.585 94.910 ;
        RECT 303.380 94.480 304.610 94.650 ;
        RECT 302.170 93.760 303.180 93.930 ;
        RECT 303.350 93.915 304.100 94.105 ;
        RECT 301.830 93.420 302.955 93.590 ;
        RECT 303.350 93.250 303.520 93.915 ;
        RECT 304.270 93.670 304.610 94.480 ;
        RECT 304.780 94.190 305.135 94.560 ;
        RECT 305.415 94.550 305.585 94.740 ;
        RECT 305.755 94.715 306.010 95.290 ;
        RECT 305.415 94.220 305.670 94.550 ;
        RECT 305.415 94.010 305.585 94.220 ;
        RECT 301.490 93.080 303.520 93.250 ;
        RECT 303.690 92.910 303.860 93.670 ;
        RECT 304.095 93.260 304.610 93.670 ;
        RECT 304.870 93.840 305.585 94.010 ;
        RECT 305.840 93.985 306.010 94.715 ;
        RECT 306.185 94.620 306.445 95.460 ;
        RECT 307.170 94.910 307.340 95.290 ;
        RECT 307.555 95.080 307.885 95.460 ;
        RECT 307.170 94.740 307.885 94.910 ;
        RECT 307.080 94.190 307.435 94.560 ;
        RECT 307.715 94.550 307.885 94.740 ;
        RECT 308.055 94.715 308.310 95.290 ;
        RECT 307.715 94.220 307.970 94.550 ;
        RECT 304.870 93.080 305.040 93.840 ;
        RECT 305.255 92.910 305.585 93.670 ;
        RECT 305.755 93.080 306.010 93.985 ;
        RECT 306.185 92.910 306.445 94.060 ;
        RECT 307.715 94.010 307.885 94.220 ;
        RECT 307.170 93.840 307.885 94.010 ;
        RECT 308.140 93.985 308.310 94.715 ;
        RECT 308.485 94.620 308.745 95.460 ;
        RECT 309.840 94.710 311.050 95.460 ;
        RECT 307.170 93.080 307.340 93.840 ;
        RECT 307.555 92.910 307.885 93.670 ;
        RECT 308.055 93.080 308.310 93.985 ;
        RECT 308.485 92.910 308.745 94.060 ;
        RECT 309.840 94.000 310.360 94.540 ;
        RECT 310.530 94.170 311.050 94.710 ;
        RECT 309.840 92.910 311.050 94.000 ;
        RECT 162.095 92.740 311.135 92.910 ;
        RECT 162.180 91.650 163.390 92.740 ;
        RECT 163.560 92.305 168.905 92.740 ;
        RECT 162.180 90.940 162.700 91.480 ;
        RECT 162.870 91.110 163.390 91.650 ;
        RECT 162.180 90.190 163.390 90.940 ;
        RECT 165.145 90.735 165.485 91.565 ;
        RECT 166.965 91.055 167.315 92.305 ;
        RECT 169.080 91.650 170.750 92.740 ;
        RECT 169.080 90.960 169.830 91.480 ;
        RECT 170.000 91.130 170.750 91.650 ;
        RECT 170.925 91.600 171.260 92.570 ;
        RECT 171.430 91.600 171.600 92.740 ;
        RECT 171.770 92.400 173.800 92.570 ;
        RECT 163.560 90.190 168.905 90.735 ;
        RECT 169.080 90.190 170.750 90.960 ;
        RECT 170.925 90.930 171.095 91.600 ;
        RECT 171.770 91.430 171.940 92.400 ;
        RECT 171.265 91.100 171.520 91.430 ;
        RECT 171.745 91.100 171.940 91.430 ;
        RECT 172.110 92.060 173.235 92.230 ;
        RECT 171.350 90.930 171.520 91.100 ;
        RECT 172.110 90.930 172.280 92.060 ;
        RECT 170.925 90.360 171.180 90.930 ;
        RECT 171.350 90.760 172.280 90.930 ;
        RECT 172.450 91.720 173.460 91.890 ;
        RECT 172.450 90.920 172.620 91.720 ;
        RECT 172.825 91.040 173.100 91.520 ;
        RECT 172.820 90.870 173.100 91.040 ;
        RECT 172.105 90.725 172.280 90.760 ;
        RECT 171.350 90.190 171.680 90.590 ;
        RECT 172.105 90.360 172.635 90.725 ;
        RECT 172.825 90.360 173.100 90.870 ;
        RECT 173.270 90.360 173.460 91.720 ;
        RECT 173.630 91.735 173.800 92.400 ;
        RECT 173.970 91.980 174.140 92.740 ;
        RECT 174.375 91.980 174.890 92.390 ;
        RECT 173.630 91.545 174.380 91.735 ;
        RECT 174.550 91.170 174.890 91.980 ;
        RECT 175.060 91.575 175.350 92.740 ;
        RECT 175.525 91.600 175.860 92.570 ;
        RECT 176.030 91.600 176.200 92.740 ;
        RECT 176.370 92.400 178.400 92.570 ;
        RECT 173.660 91.000 174.890 91.170 ;
        RECT 173.640 90.190 174.150 90.725 ;
        RECT 174.370 90.395 174.615 91.000 ;
        RECT 175.525 90.930 175.695 91.600 ;
        RECT 176.370 91.430 176.540 92.400 ;
        RECT 175.865 91.100 176.120 91.430 ;
        RECT 176.345 91.100 176.540 91.430 ;
        RECT 176.710 92.060 177.835 92.230 ;
        RECT 175.950 90.930 176.120 91.100 ;
        RECT 176.710 90.930 176.880 92.060 ;
        RECT 175.060 90.190 175.350 90.915 ;
        RECT 175.525 90.360 175.780 90.930 ;
        RECT 175.950 90.760 176.880 90.930 ;
        RECT 177.050 91.720 178.060 91.890 ;
        RECT 177.050 90.920 177.220 91.720 ;
        RECT 177.425 91.040 177.700 91.520 ;
        RECT 177.420 90.870 177.700 91.040 ;
        RECT 176.705 90.725 176.880 90.760 ;
        RECT 175.950 90.190 176.280 90.590 ;
        RECT 176.705 90.360 177.235 90.725 ;
        RECT 177.425 90.360 177.700 90.870 ;
        RECT 177.870 90.360 178.060 91.720 ;
        RECT 178.230 91.735 178.400 92.400 ;
        RECT 178.570 91.980 178.740 92.740 ;
        RECT 178.975 91.980 179.490 92.390 ;
        RECT 178.230 91.545 178.980 91.735 ;
        RECT 179.150 91.170 179.490 91.980 ;
        RECT 178.260 91.000 179.490 91.170 ;
        RECT 179.660 91.600 180.045 92.570 ;
        RECT 180.215 92.280 180.540 92.740 ;
        RECT 181.060 92.110 181.340 92.570 ;
        RECT 180.215 91.890 181.340 92.110 ;
        RECT 178.240 90.190 178.750 90.725 ;
        RECT 178.970 90.395 179.215 91.000 ;
        RECT 179.660 90.930 179.940 91.600 ;
        RECT 180.215 91.430 180.665 91.890 ;
        RECT 181.530 91.720 181.930 92.570 ;
        RECT 182.330 92.280 182.600 92.740 ;
        RECT 182.770 92.110 183.055 92.570 ;
        RECT 180.110 91.100 180.665 91.430 ;
        RECT 180.835 91.160 181.930 91.720 ;
        RECT 180.215 90.990 180.665 91.100 ;
        RECT 179.660 90.360 180.045 90.930 ;
        RECT 180.215 90.820 181.340 90.990 ;
        RECT 180.215 90.190 180.540 90.650 ;
        RECT 181.060 90.360 181.340 90.820 ;
        RECT 181.530 90.360 181.930 91.160 ;
        RECT 182.100 91.890 183.055 92.110 ;
        RECT 183.345 92.070 183.600 92.570 ;
        RECT 183.770 92.240 184.100 92.740 ;
        RECT 183.345 91.900 184.095 92.070 ;
        RECT 182.100 90.990 182.310 91.890 ;
        RECT 182.480 91.160 183.170 91.720 ;
        RECT 183.345 91.080 183.695 91.730 ;
        RECT 182.100 90.820 183.055 90.990 ;
        RECT 183.865 90.910 184.095 91.900 ;
        RECT 182.330 90.190 182.600 90.650 ;
        RECT 182.770 90.360 183.055 90.820 ;
        RECT 183.345 90.740 184.095 90.910 ;
        RECT 183.345 90.450 183.600 90.740 ;
        RECT 183.770 90.190 184.100 90.570 ;
        RECT 184.270 90.450 184.440 92.570 ;
        RECT 184.610 91.770 184.935 92.555 ;
        RECT 185.105 92.280 185.355 92.740 ;
        RECT 185.525 92.240 185.775 92.570 ;
        RECT 185.990 92.240 186.670 92.570 ;
        RECT 185.525 92.110 185.695 92.240 ;
        RECT 185.300 91.940 185.695 92.110 ;
        RECT 184.670 90.720 185.130 91.770 ;
        RECT 185.300 90.580 185.470 91.940 ;
        RECT 185.865 91.680 186.330 92.070 ;
        RECT 185.640 90.870 185.990 91.490 ;
        RECT 186.160 91.090 186.330 91.680 ;
        RECT 186.500 91.460 186.670 92.240 ;
        RECT 186.840 92.140 187.010 92.480 ;
        RECT 187.245 92.310 187.575 92.740 ;
        RECT 187.745 92.140 187.915 92.480 ;
        RECT 188.210 92.280 188.580 92.740 ;
        RECT 186.840 91.970 187.915 92.140 ;
        RECT 188.750 92.110 188.920 92.570 ;
        RECT 189.155 92.230 190.025 92.570 ;
        RECT 190.195 92.280 190.445 92.740 ;
        RECT 188.360 91.940 188.920 92.110 ;
        RECT 188.360 91.800 188.530 91.940 ;
        RECT 187.030 91.630 188.530 91.800 ;
        RECT 189.225 91.770 189.685 92.060 ;
        RECT 186.500 91.290 188.190 91.460 ;
        RECT 186.160 90.870 186.515 91.090 ;
        RECT 186.685 90.580 186.855 91.290 ;
        RECT 187.060 90.870 187.850 91.120 ;
        RECT 188.020 91.110 188.190 91.290 ;
        RECT 188.360 90.940 188.530 91.630 ;
        RECT 184.800 90.190 185.130 90.550 ;
        RECT 185.300 90.410 185.795 90.580 ;
        RECT 186.000 90.410 186.855 90.580 ;
        RECT 187.730 90.190 188.060 90.650 ;
        RECT 188.270 90.550 188.530 90.940 ;
        RECT 188.720 91.760 189.685 91.770 ;
        RECT 189.855 91.850 190.025 92.230 ;
        RECT 190.615 92.190 190.785 92.480 ;
        RECT 190.965 92.360 191.295 92.740 ;
        RECT 190.615 92.020 191.415 92.190 ;
        RECT 188.720 91.600 189.395 91.760 ;
        RECT 189.855 91.680 191.075 91.850 ;
        RECT 188.720 90.810 188.930 91.600 ;
        RECT 189.855 91.590 190.025 91.680 ;
        RECT 189.100 90.810 189.450 91.430 ;
        RECT 189.620 91.420 190.025 91.590 ;
        RECT 189.620 90.640 189.790 91.420 ;
        RECT 189.960 90.970 190.180 91.250 ;
        RECT 190.360 91.140 190.900 91.510 ;
        RECT 191.245 91.430 191.415 92.020 ;
        RECT 191.635 91.600 191.940 92.740 ;
        RECT 192.110 91.550 192.365 92.430 ;
        RECT 192.540 91.650 194.210 92.740 ;
        RECT 191.245 91.400 191.985 91.430 ;
        RECT 189.960 90.800 190.490 90.970 ;
        RECT 188.270 90.380 188.620 90.550 ;
        RECT 188.840 90.360 189.790 90.640 ;
        RECT 189.960 90.190 190.150 90.630 ;
        RECT 190.320 90.570 190.490 90.800 ;
        RECT 190.660 90.740 190.900 91.140 ;
        RECT 191.070 91.100 191.985 91.400 ;
        RECT 191.070 90.925 191.395 91.100 ;
        RECT 191.070 90.570 191.390 90.925 ;
        RECT 192.155 90.900 192.365 91.550 ;
        RECT 190.320 90.400 191.390 90.570 ;
        RECT 191.635 90.190 191.940 90.650 ;
        RECT 192.110 90.370 192.365 90.900 ;
        RECT 192.540 90.960 193.290 91.480 ;
        RECT 193.460 91.130 194.210 91.650 ;
        RECT 195.045 91.770 195.375 92.570 ;
        RECT 195.545 91.940 195.875 92.740 ;
        RECT 196.175 91.770 196.505 92.570 ;
        RECT 197.150 91.940 197.400 92.740 ;
        RECT 195.045 91.600 197.480 91.770 ;
        RECT 197.670 91.600 197.840 92.740 ;
        RECT 198.010 91.600 198.350 92.570 ;
        RECT 198.520 91.650 200.190 92.740 ;
        RECT 194.840 91.180 195.190 91.430 ;
        RECT 195.375 90.970 195.545 91.600 ;
        RECT 195.715 91.180 196.045 91.380 ;
        RECT 196.215 91.180 196.545 91.380 ;
        RECT 196.715 91.180 197.135 91.380 ;
        RECT 197.310 91.350 197.480 91.600 ;
        RECT 197.310 91.180 198.005 91.350 ;
        RECT 192.540 90.190 194.210 90.960 ;
        RECT 195.045 90.360 195.545 90.970 ;
        RECT 196.175 90.840 197.400 91.010 ;
        RECT 198.175 90.990 198.350 91.600 ;
        RECT 196.175 90.360 196.505 90.840 ;
        RECT 196.675 90.190 196.900 90.650 ;
        RECT 197.070 90.360 197.400 90.840 ;
        RECT 197.590 90.190 197.840 90.990 ;
        RECT 198.010 90.360 198.350 90.990 ;
        RECT 198.520 90.960 199.270 91.480 ;
        RECT 199.440 91.130 200.190 91.650 ;
        RECT 200.820 91.575 201.110 92.740 ;
        RECT 201.280 91.650 203.870 92.740 ;
        RECT 201.280 90.960 202.490 91.480 ;
        RECT 202.660 91.130 203.870 91.650 ;
        RECT 204.130 91.810 204.300 92.570 ;
        RECT 204.515 91.980 204.845 92.740 ;
        RECT 204.130 91.640 204.845 91.810 ;
        RECT 205.015 91.665 205.270 92.570 ;
        RECT 204.040 91.090 204.395 91.460 ;
        RECT 204.675 91.430 204.845 91.640 ;
        RECT 204.675 91.100 204.930 91.430 ;
        RECT 198.520 90.190 200.190 90.960 ;
        RECT 200.820 90.190 201.110 90.915 ;
        RECT 201.280 90.190 203.870 90.960 ;
        RECT 204.675 90.910 204.845 91.100 ;
        RECT 205.100 90.935 205.270 91.665 ;
        RECT 205.445 91.590 205.705 92.740 ;
        RECT 206.360 91.850 206.620 92.560 ;
        RECT 206.790 92.030 207.120 92.740 ;
        RECT 207.290 91.850 207.520 92.560 ;
        RECT 206.360 91.610 207.520 91.850 ;
        RECT 207.700 91.830 207.970 92.560 ;
        RECT 208.150 92.010 208.490 92.740 ;
        RECT 207.700 91.610 208.470 91.830 ;
        RECT 206.350 91.100 206.650 91.430 ;
        RECT 206.830 91.120 207.355 91.430 ;
        RECT 207.535 91.120 208.000 91.430 ;
        RECT 204.130 90.740 204.845 90.910 ;
        RECT 204.130 90.360 204.300 90.740 ;
        RECT 204.515 90.190 204.845 90.570 ;
        RECT 205.015 90.360 205.270 90.935 ;
        RECT 205.445 90.190 205.705 91.030 ;
        RECT 206.360 90.190 206.650 90.920 ;
        RECT 206.830 90.480 207.060 91.120 ;
        RECT 208.180 90.940 208.470 91.610 ;
        RECT 207.240 90.740 208.470 90.940 ;
        RECT 207.240 90.370 207.550 90.740 ;
        RECT 207.730 90.190 208.400 90.560 ;
        RECT 208.660 90.370 208.920 92.560 ;
        RECT 209.255 91.730 209.555 92.570 ;
        RECT 209.750 91.900 210.000 92.740 ;
        RECT 210.590 92.150 211.395 92.570 ;
        RECT 210.170 91.980 211.735 92.150 ;
        RECT 210.170 91.730 210.340 91.980 ;
        RECT 209.255 91.560 210.340 91.730 ;
        RECT 209.100 91.100 209.430 91.390 ;
        RECT 209.600 90.930 209.770 91.560 ;
        RECT 210.510 91.430 210.830 91.810 ;
        RECT 209.940 91.180 210.270 91.390 ;
        RECT 210.450 91.180 210.830 91.430 ;
        RECT 211.020 91.390 211.395 91.810 ;
        RECT 211.565 91.730 211.735 91.980 ;
        RECT 211.905 91.900 212.235 92.740 ;
        RECT 212.405 91.980 213.070 92.570 ;
        RECT 213.240 92.305 218.585 92.740 ;
        RECT 211.565 91.560 212.485 91.730 ;
        RECT 212.315 91.390 212.485 91.560 ;
        RECT 211.020 91.380 211.505 91.390 ;
        RECT 211.000 91.210 211.505 91.380 ;
        RECT 211.020 91.180 211.505 91.210 ;
        RECT 211.695 91.180 212.145 91.390 ;
        RECT 212.315 91.180 212.650 91.390 ;
        RECT 212.820 91.010 213.070 91.980 ;
        RECT 209.260 90.750 209.770 90.930 ;
        RECT 210.175 90.840 211.875 91.010 ;
        RECT 210.175 90.750 210.560 90.840 ;
        RECT 209.260 90.360 209.590 90.750 ;
        RECT 209.760 90.410 210.945 90.580 ;
        RECT 211.205 90.190 211.375 90.660 ;
        RECT 211.545 90.375 211.875 90.840 ;
        RECT 212.045 90.190 212.215 91.010 ;
        RECT 212.385 90.370 213.070 91.010 ;
        RECT 214.825 90.735 215.165 91.565 ;
        RECT 216.645 91.055 216.995 92.305 ;
        RECT 218.760 91.650 222.270 92.740 ;
        RECT 218.760 90.960 220.410 91.480 ;
        RECT 220.580 91.130 222.270 91.650 ;
        RECT 223.360 91.890 223.620 92.570 ;
        RECT 223.790 91.960 224.040 92.740 ;
        RECT 224.290 92.190 224.540 92.570 ;
        RECT 224.710 92.360 225.065 92.740 ;
        RECT 226.070 92.350 226.405 92.570 ;
        RECT 225.670 92.190 225.900 92.230 ;
        RECT 224.290 91.990 225.900 92.190 ;
        RECT 224.290 91.980 225.125 91.990 ;
        RECT 225.715 91.900 225.900 91.990 ;
        RECT 213.240 90.190 218.585 90.735 ;
        RECT 218.760 90.190 222.270 90.960 ;
        RECT 223.360 90.700 223.530 91.890 ;
        RECT 225.230 91.790 225.560 91.820 ;
        RECT 223.760 91.730 225.560 91.790 ;
        RECT 226.150 91.730 226.405 92.350 ;
        RECT 223.700 91.620 226.405 91.730 ;
        RECT 223.700 91.585 223.900 91.620 ;
        RECT 223.700 91.010 223.870 91.585 ;
        RECT 225.230 91.560 226.405 91.620 ;
        RECT 226.580 91.575 226.870 92.740 ;
        RECT 227.060 91.900 227.315 92.570 ;
        RECT 227.485 91.980 227.815 92.740 ;
        RECT 227.985 92.140 228.235 92.570 ;
        RECT 228.405 92.320 228.760 92.740 ;
        RECT 228.950 92.400 230.120 92.570 ;
        RECT 228.950 92.360 229.280 92.400 ;
        RECT 229.390 92.140 229.620 92.230 ;
        RECT 227.985 91.900 229.620 92.140 ;
        RECT 229.790 91.900 230.120 92.400 ;
        RECT 224.100 91.145 224.510 91.450 ;
        RECT 224.680 91.180 225.010 91.390 ;
        RECT 223.700 90.890 223.970 91.010 ;
        RECT 223.700 90.845 224.545 90.890 ;
        RECT 223.790 90.720 224.545 90.845 ;
        RECT 224.800 90.780 225.010 91.180 ;
        RECT 225.255 91.180 225.730 91.390 ;
        RECT 225.920 91.180 226.410 91.380 ;
        RECT 225.255 90.780 225.475 91.180 ;
        RECT 223.360 90.690 223.590 90.700 ;
        RECT 223.360 90.360 223.620 90.690 ;
        RECT 224.375 90.570 224.545 90.720 ;
        RECT 223.790 90.190 224.120 90.550 ;
        RECT 224.375 90.360 225.675 90.570 ;
        RECT 225.950 90.190 226.405 90.955 ;
        RECT 226.580 90.190 226.870 90.915 ;
        RECT 227.060 90.770 227.230 91.900 ;
        RECT 230.290 91.730 230.460 92.570 ;
        RECT 227.400 91.560 230.460 91.730 ;
        RECT 230.720 91.890 230.980 92.570 ;
        RECT 231.150 91.960 231.400 92.740 ;
        RECT 231.650 92.190 231.900 92.570 ;
        RECT 232.070 92.360 232.425 92.740 ;
        RECT 233.430 92.350 233.765 92.570 ;
        RECT 233.030 92.190 233.260 92.230 ;
        RECT 231.650 91.990 233.260 92.190 ;
        RECT 231.650 91.980 232.485 91.990 ;
        RECT 233.075 91.900 233.260 91.990 ;
        RECT 227.400 91.010 227.570 91.560 ;
        RECT 227.800 91.180 228.165 91.380 ;
        RECT 228.335 91.180 228.665 91.380 ;
        RECT 227.400 90.840 228.200 91.010 ;
        RECT 227.060 90.700 227.245 90.770 ;
        RECT 227.060 90.690 227.270 90.700 ;
        RECT 227.060 90.360 227.315 90.690 ;
        RECT 227.530 90.190 227.860 90.670 ;
        RECT 228.030 90.610 228.200 90.840 ;
        RECT 228.380 90.780 228.665 91.180 ;
        RECT 228.935 91.180 229.410 91.380 ;
        RECT 229.580 91.180 230.025 91.380 ;
        RECT 230.195 91.180 230.545 91.390 ;
        RECT 228.935 90.780 229.215 91.180 ;
        RECT 229.395 90.840 230.460 91.010 ;
        RECT 229.395 90.610 229.565 90.840 ;
        RECT 228.030 90.360 229.565 90.610 ;
        RECT 229.790 90.190 230.120 90.670 ;
        RECT 230.290 90.360 230.460 90.840 ;
        RECT 230.720 90.700 230.890 91.890 ;
        RECT 232.590 91.790 232.920 91.820 ;
        RECT 231.120 91.730 232.920 91.790 ;
        RECT 233.510 91.730 233.765 92.350 ;
        RECT 233.940 92.305 239.285 92.740 ;
        RECT 231.060 91.620 233.765 91.730 ;
        RECT 231.060 91.585 231.260 91.620 ;
        RECT 231.060 91.010 231.230 91.585 ;
        RECT 232.590 91.560 233.765 91.620 ;
        RECT 231.460 91.145 231.870 91.450 ;
        RECT 232.040 91.180 232.370 91.390 ;
        RECT 231.060 90.890 231.330 91.010 ;
        RECT 231.060 90.845 231.905 90.890 ;
        RECT 231.150 90.720 231.905 90.845 ;
        RECT 232.160 90.780 232.370 91.180 ;
        RECT 232.615 91.180 233.090 91.390 ;
        RECT 233.280 91.180 233.770 91.380 ;
        RECT 232.615 90.780 232.835 91.180 ;
        RECT 230.720 90.690 230.950 90.700 ;
        RECT 230.720 90.360 230.980 90.690 ;
        RECT 231.735 90.570 231.905 90.720 ;
        RECT 231.150 90.190 231.480 90.550 ;
        RECT 231.735 90.360 233.035 90.570 ;
        RECT 233.310 90.190 233.765 90.955 ;
        RECT 235.525 90.735 235.865 91.565 ;
        RECT 237.345 91.055 237.695 92.305 ;
        RECT 239.460 91.650 241.130 92.740 ;
        RECT 239.460 90.960 240.210 91.480 ;
        RECT 240.380 91.130 241.130 91.650 ;
        RECT 241.305 92.020 241.640 92.530 ;
        RECT 233.940 90.190 239.285 90.735 ;
        RECT 239.460 90.190 241.130 90.960 ;
        RECT 241.305 90.665 241.560 92.020 ;
        RECT 241.890 91.940 242.220 92.740 ;
        RECT 242.465 92.150 242.750 92.570 ;
        RECT 243.005 92.320 243.335 92.740 ;
        RECT 243.560 92.400 244.720 92.570 ;
        RECT 243.560 92.150 243.890 92.400 ;
        RECT 242.465 91.980 243.890 92.150 ;
        RECT 244.120 91.770 244.290 92.230 ;
        RECT 244.550 91.900 244.720 92.400 ;
        RECT 245.000 91.900 245.255 92.570 ;
        RECT 245.425 91.980 245.755 92.740 ;
        RECT 245.925 92.140 246.175 92.570 ;
        RECT 246.345 92.320 246.700 92.740 ;
        RECT 246.890 92.400 248.060 92.570 ;
        RECT 246.890 92.360 247.220 92.400 ;
        RECT 247.330 92.140 247.560 92.230 ;
        RECT 245.925 91.900 247.560 92.140 ;
        RECT 247.730 91.900 248.060 92.400 ;
        RECT 241.920 91.600 244.290 91.770 ;
        RECT 245.000 91.890 245.210 91.900 ;
        RECT 241.920 91.430 242.090 91.600 ;
        RECT 244.540 91.430 244.745 91.720 ;
        RECT 241.785 91.100 242.090 91.430 ;
        RECT 242.285 91.380 242.535 91.430 ;
        RECT 242.745 91.380 243.015 91.430 ;
        RECT 242.280 91.210 242.535 91.380 ;
        RECT 242.740 91.210 243.015 91.380 ;
        RECT 242.285 91.100 242.535 91.210 ;
        RECT 241.920 90.930 242.090 91.100 ;
        RECT 241.920 90.760 242.480 90.930 ;
        RECT 242.745 90.770 243.015 91.210 ;
        RECT 243.205 91.040 243.495 91.430 ;
        RECT 243.200 90.870 243.495 91.040 ;
        RECT 243.205 90.770 243.495 90.870 ;
        RECT 243.665 90.765 244.085 91.430 ;
        RECT 244.395 91.380 244.745 91.430 ;
        RECT 244.395 91.210 244.750 91.380 ;
        RECT 244.395 91.100 244.745 91.210 ;
        RECT 241.305 90.405 241.640 90.665 ;
        RECT 242.310 90.590 242.480 90.760 ;
        RECT 241.810 90.190 242.140 90.590 ;
        RECT 242.310 90.420 243.925 90.590 ;
        RECT 244.470 90.190 244.800 90.910 ;
        RECT 245.000 90.770 245.170 91.890 ;
        RECT 248.230 91.730 248.400 92.570 ;
        RECT 245.340 91.560 248.400 91.730 ;
        RECT 248.660 91.650 252.170 92.740 ;
        RECT 245.340 91.010 245.510 91.560 ;
        RECT 245.740 91.180 246.105 91.380 ;
        RECT 246.275 91.180 246.605 91.380 ;
        RECT 245.340 90.840 246.140 91.010 ;
        RECT 245.000 90.690 245.185 90.770 ;
        RECT 245.000 90.360 245.255 90.690 ;
        RECT 245.470 90.190 245.800 90.670 ;
        RECT 245.970 90.610 246.140 90.840 ;
        RECT 246.320 90.780 246.605 91.180 ;
        RECT 246.875 91.180 247.350 91.380 ;
        RECT 247.520 91.180 247.965 91.380 ;
        RECT 248.135 91.180 248.485 91.390 ;
        RECT 246.875 90.780 247.155 91.180 ;
        RECT 247.335 90.840 248.400 91.010 ;
        RECT 247.335 90.610 247.505 90.840 ;
        RECT 245.970 90.360 247.505 90.610 ;
        RECT 247.730 90.190 248.060 90.670 ;
        RECT 248.230 90.360 248.400 90.840 ;
        RECT 248.660 90.960 250.310 91.480 ;
        RECT 250.480 91.130 252.170 91.650 ;
        RECT 252.340 91.575 252.630 92.740 ;
        RECT 252.800 92.305 258.145 92.740 ;
        RECT 248.660 90.190 252.170 90.960 ;
        RECT 252.340 90.190 252.630 90.915 ;
        RECT 254.385 90.735 254.725 91.565 ;
        RECT 256.205 91.055 256.555 92.305 ;
        RECT 258.870 91.730 259.040 92.570 ;
        RECT 259.210 92.400 260.380 92.570 ;
        RECT 259.210 91.900 259.540 92.400 ;
        RECT 260.050 92.360 260.380 92.400 ;
        RECT 260.570 92.320 260.925 92.740 ;
        RECT 259.710 92.140 259.940 92.230 ;
        RECT 261.095 92.140 261.345 92.570 ;
        RECT 259.710 91.900 261.345 92.140 ;
        RECT 261.515 91.980 261.845 92.740 ;
        RECT 262.015 91.900 262.270 92.570 ;
        RECT 258.870 91.560 261.930 91.730 ;
        RECT 258.785 91.180 259.135 91.390 ;
        RECT 259.305 91.180 259.750 91.380 ;
        RECT 259.920 91.180 260.395 91.380 ;
        RECT 258.870 90.840 259.935 91.010 ;
        RECT 252.800 90.190 258.145 90.735 ;
        RECT 258.870 90.360 259.040 90.840 ;
        RECT 259.210 90.190 259.540 90.670 ;
        RECT 259.765 90.610 259.935 90.840 ;
        RECT 260.115 90.780 260.395 91.180 ;
        RECT 260.665 91.180 260.995 91.380 ;
        RECT 261.165 91.180 261.530 91.380 ;
        RECT 260.665 90.780 260.950 91.180 ;
        RECT 261.760 91.010 261.930 91.560 ;
        RECT 261.130 90.840 261.930 91.010 ;
        RECT 261.130 90.610 261.300 90.840 ;
        RECT 262.100 90.770 262.270 91.900 ;
        RECT 262.465 92.350 262.800 92.570 ;
        RECT 263.805 92.360 264.160 92.740 ;
        RECT 262.465 91.730 262.720 92.350 ;
        RECT 262.970 92.190 263.200 92.230 ;
        RECT 264.330 92.190 264.580 92.570 ;
        RECT 262.970 91.990 264.580 92.190 ;
        RECT 262.970 91.900 263.155 91.990 ;
        RECT 263.745 91.980 264.580 91.990 ;
        RECT 264.830 91.960 265.080 92.740 ;
        RECT 265.250 91.890 265.510 92.570 ;
        RECT 263.310 91.790 263.640 91.820 ;
        RECT 263.310 91.730 265.110 91.790 ;
        RECT 262.465 91.620 265.170 91.730 ;
        RECT 262.465 91.560 263.640 91.620 ;
        RECT 264.970 91.585 265.170 91.620 ;
        RECT 262.460 91.180 262.950 91.380 ;
        RECT 263.140 91.180 263.615 91.390 ;
        RECT 262.085 90.690 262.270 90.770 ;
        RECT 259.765 90.360 261.300 90.610 ;
        RECT 261.470 90.190 261.800 90.670 ;
        RECT 262.015 90.360 262.270 90.690 ;
        RECT 262.465 90.190 262.920 90.955 ;
        RECT 263.395 90.780 263.615 91.180 ;
        RECT 263.860 91.180 264.190 91.390 ;
        RECT 263.860 90.780 264.070 91.180 ;
        RECT 264.360 91.145 264.770 91.450 ;
        RECT 265.000 91.010 265.170 91.585 ;
        RECT 264.900 90.890 265.170 91.010 ;
        RECT 264.325 90.845 265.170 90.890 ;
        RECT 264.325 90.720 265.080 90.845 ;
        RECT 264.325 90.570 264.495 90.720 ;
        RECT 265.340 90.700 265.510 91.890 ;
        RECT 265.685 92.350 266.020 92.570 ;
        RECT 267.025 92.360 267.380 92.740 ;
        RECT 265.685 91.730 265.940 92.350 ;
        RECT 266.190 92.190 266.420 92.230 ;
        RECT 267.550 92.190 267.800 92.570 ;
        RECT 266.190 91.990 267.800 92.190 ;
        RECT 266.190 91.900 266.375 91.990 ;
        RECT 266.965 91.980 267.800 91.990 ;
        RECT 268.050 91.960 268.300 92.740 ;
        RECT 268.470 91.890 268.730 92.570 ;
        RECT 268.900 92.305 274.245 92.740 ;
        RECT 266.530 91.790 266.860 91.820 ;
        RECT 266.530 91.730 268.330 91.790 ;
        RECT 265.685 91.620 268.390 91.730 ;
        RECT 265.685 91.560 266.860 91.620 ;
        RECT 268.190 91.585 268.390 91.620 ;
        RECT 265.680 91.180 266.170 91.380 ;
        RECT 266.360 91.180 266.835 91.390 ;
        RECT 265.280 90.690 265.510 90.700 ;
        RECT 263.195 90.360 264.495 90.570 ;
        RECT 264.750 90.190 265.080 90.550 ;
        RECT 265.250 90.360 265.510 90.690 ;
        RECT 265.685 90.190 266.140 90.955 ;
        RECT 266.615 90.780 266.835 91.180 ;
        RECT 267.080 91.180 267.410 91.390 ;
        RECT 267.080 90.780 267.290 91.180 ;
        RECT 267.580 91.145 267.990 91.450 ;
        RECT 268.220 91.010 268.390 91.585 ;
        RECT 268.120 90.890 268.390 91.010 ;
        RECT 267.545 90.845 268.390 90.890 ;
        RECT 267.545 90.720 268.300 90.845 ;
        RECT 267.545 90.570 267.715 90.720 ;
        RECT 268.560 90.700 268.730 91.890 ;
        RECT 270.485 90.735 270.825 91.565 ;
        RECT 272.305 91.055 272.655 92.305 ;
        RECT 274.420 91.650 277.930 92.740 ;
        RECT 274.420 90.960 276.070 91.480 ;
        RECT 276.240 91.130 277.930 91.650 ;
        RECT 278.100 91.575 278.390 92.740 ;
        RECT 278.565 92.020 278.900 92.530 ;
        RECT 268.500 90.690 268.730 90.700 ;
        RECT 266.415 90.360 267.715 90.570 ;
        RECT 267.970 90.190 268.300 90.550 ;
        RECT 268.470 90.360 268.730 90.690 ;
        RECT 268.900 90.190 274.245 90.735 ;
        RECT 274.420 90.190 277.930 90.960 ;
        RECT 278.100 90.190 278.390 90.915 ;
        RECT 278.565 90.665 278.820 92.020 ;
        RECT 279.150 91.940 279.480 92.740 ;
        RECT 279.725 92.150 280.010 92.570 ;
        RECT 280.265 92.320 280.595 92.740 ;
        RECT 280.820 92.400 281.980 92.570 ;
        RECT 280.820 92.150 281.150 92.400 ;
        RECT 279.725 91.980 281.150 92.150 ;
        RECT 281.380 91.770 281.550 92.230 ;
        RECT 281.810 91.900 281.980 92.400 ;
        RECT 279.180 91.600 281.550 91.770 ;
        RECT 279.180 91.430 279.350 91.600 ;
        RECT 281.800 91.550 282.010 91.720 ;
        RECT 282.240 91.650 285.750 92.740 ;
        RECT 281.800 91.430 282.005 91.550 ;
        RECT 279.045 91.100 279.350 91.430 ;
        RECT 279.545 91.380 279.795 91.430 ;
        RECT 280.005 91.380 280.275 91.430 ;
        RECT 279.540 91.210 279.795 91.380 ;
        RECT 280.000 91.210 280.275 91.380 ;
        RECT 279.545 91.100 279.795 91.210 ;
        RECT 279.180 90.930 279.350 91.100 ;
        RECT 279.180 90.760 279.740 90.930 ;
        RECT 280.005 90.770 280.275 91.210 ;
        RECT 280.465 91.040 280.755 91.430 ;
        RECT 280.460 90.870 280.755 91.040 ;
        RECT 280.465 90.770 280.755 90.870 ;
        RECT 280.925 90.765 281.345 91.430 ;
        RECT 281.655 91.100 282.005 91.430 ;
        RECT 282.240 90.960 283.890 91.480 ;
        RECT 284.060 91.130 285.750 91.650 ;
        RECT 286.385 91.550 286.640 92.430 ;
        RECT 286.810 91.600 287.115 92.740 ;
        RECT 287.455 92.360 287.785 92.740 ;
        RECT 287.965 92.190 288.135 92.480 ;
        RECT 288.305 92.280 288.555 92.740 ;
        RECT 287.335 92.020 288.135 92.190 ;
        RECT 288.725 92.230 289.595 92.570 ;
        RECT 278.565 90.405 278.900 90.665 ;
        RECT 279.570 90.590 279.740 90.760 ;
        RECT 279.070 90.190 279.400 90.590 ;
        RECT 279.570 90.420 281.185 90.590 ;
        RECT 281.730 90.190 282.060 90.910 ;
        RECT 282.240 90.190 285.750 90.960 ;
        RECT 286.385 90.900 286.595 91.550 ;
        RECT 287.335 91.430 287.505 92.020 ;
        RECT 288.725 91.850 288.895 92.230 ;
        RECT 289.830 92.110 290.000 92.570 ;
        RECT 290.170 92.280 290.540 92.740 ;
        RECT 290.835 92.140 291.005 92.480 ;
        RECT 291.175 92.310 291.505 92.740 ;
        RECT 291.740 92.140 291.910 92.480 ;
        RECT 287.675 91.680 288.895 91.850 ;
        RECT 289.065 91.770 289.525 92.060 ;
        RECT 289.830 91.940 290.390 92.110 ;
        RECT 290.835 91.970 291.910 92.140 ;
        RECT 292.080 92.240 292.760 92.570 ;
        RECT 292.975 92.240 293.225 92.570 ;
        RECT 293.395 92.280 293.645 92.740 ;
        RECT 290.220 91.800 290.390 91.940 ;
        RECT 289.065 91.760 290.030 91.770 ;
        RECT 288.725 91.590 288.895 91.680 ;
        RECT 289.355 91.600 290.030 91.760 ;
        RECT 286.765 91.400 287.505 91.430 ;
        RECT 286.765 91.100 287.680 91.400 ;
        RECT 287.355 90.925 287.680 91.100 ;
        RECT 286.385 90.370 286.640 90.900 ;
        RECT 286.810 90.190 287.115 90.650 ;
        RECT 287.360 90.570 287.680 90.925 ;
        RECT 287.850 91.140 288.390 91.510 ;
        RECT 288.725 91.420 289.130 91.590 ;
        RECT 287.850 90.740 288.090 91.140 ;
        RECT 288.570 90.970 288.790 91.250 ;
        RECT 288.260 90.800 288.790 90.970 ;
        RECT 288.260 90.570 288.430 90.800 ;
        RECT 288.960 90.640 289.130 91.420 ;
        RECT 289.300 90.810 289.650 91.430 ;
        RECT 289.820 90.810 290.030 91.600 ;
        RECT 290.220 91.630 291.720 91.800 ;
        RECT 290.220 90.940 290.390 91.630 ;
        RECT 292.080 91.460 292.250 92.240 ;
        RECT 293.055 92.110 293.225 92.240 ;
        RECT 290.560 91.290 292.250 91.460 ;
        RECT 292.420 91.680 292.885 92.070 ;
        RECT 293.055 91.940 293.450 92.110 ;
        RECT 290.560 91.110 290.730 91.290 ;
        RECT 287.360 90.400 288.430 90.570 ;
        RECT 288.600 90.190 288.790 90.630 ;
        RECT 288.960 90.360 289.910 90.640 ;
        RECT 290.220 90.550 290.480 90.940 ;
        RECT 290.900 90.870 291.690 91.120 ;
        RECT 290.130 90.380 290.480 90.550 ;
        RECT 290.690 90.190 291.020 90.650 ;
        RECT 291.895 90.580 292.065 91.290 ;
        RECT 292.420 91.090 292.590 91.680 ;
        RECT 292.235 90.870 292.590 91.090 ;
        RECT 292.760 90.870 293.110 91.490 ;
        RECT 293.280 90.580 293.450 91.940 ;
        RECT 293.815 91.770 294.140 92.555 ;
        RECT 293.620 90.720 294.080 91.770 ;
        RECT 291.895 90.410 292.750 90.580 ;
        RECT 292.955 90.410 293.450 90.580 ;
        RECT 293.620 90.190 293.950 90.550 ;
        RECT 294.310 90.450 294.480 92.570 ;
        RECT 294.650 92.240 294.980 92.740 ;
        RECT 295.150 92.070 295.405 92.570 ;
        RECT 294.655 91.900 295.405 92.070 ;
        RECT 294.655 90.910 294.885 91.900 ;
        RECT 295.055 91.080 295.405 91.730 ;
        RECT 296.045 91.600 296.380 92.570 ;
        RECT 296.550 91.600 296.720 92.740 ;
        RECT 296.890 92.400 298.920 92.570 ;
        RECT 296.045 90.930 296.215 91.600 ;
        RECT 296.890 91.430 297.060 92.400 ;
        RECT 296.385 91.100 296.640 91.430 ;
        RECT 296.865 91.100 297.060 91.430 ;
        RECT 297.230 92.060 298.355 92.230 ;
        RECT 296.470 90.930 296.640 91.100 ;
        RECT 297.230 90.930 297.400 92.060 ;
        RECT 294.655 90.740 295.405 90.910 ;
        RECT 294.650 90.190 294.980 90.570 ;
        RECT 295.150 90.450 295.405 90.740 ;
        RECT 296.045 90.360 296.300 90.930 ;
        RECT 296.470 90.760 297.400 90.930 ;
        RECT 297.570 91.720 298.580 91.890 ;
        RECT 297.570 90.920 297.740 91.720 ;
        RECT 297.945 91.380 298.220 91.520 ;
        RECT 297.940 91.210 298.220 91.380 ;
        RECT 297.225 90.725 297.400 90.760 ;
        RECT 296.470 90.190 296.800 90.590 ;
        RECT 297.225 90.360 297.755 90.725 ;
        RECT 297.945 90.360 298.220 91.210 ;
        RECT 298.390 90.360 298.580 91.720 ;
        RECT 298.750 91.735 298.920 92.400 ;
        RECT 299.090 91.980 299.260 92.740 ;
        RECT 299.495 91.980 300.010 92.390 ;
        RECT 298.750 91.545 299.500 91.735 ;
        RECT 299.670 91.170 300.010 91.980 ;
        RECT 300.180 91.650 301.850 92.740 ;
        RECT 298.780 91.000 300.010 91.170 ;
        RECT 298.760 90.190 299.270 90.725 ;
        RECT 299.490 90.395 299.735 91.000 ;
        RECT 300.180 90.960 300.930 91.480 ;
        RECT 301.100 91.130 301.850 91.650 ;
        RECT 302.110 91.810 302.280 92.570 ;
        RECT 302.495 91.980 302.825 92.740 ;
        RECT 302.110 91.640 302.825 91.810 ;
        RECT 302.995 91.665 303.250 92.570 ;
        RECT 302.020 91.090 302.375 91.460 ;
        RECT 302.655 91.430 302.825 91.640 ;
        RECT 302.655 91.100 302.910 91.430 ;
        RECT 300.180 90.190 301.850 90.960 ;
        RECT 302.655 90.910 302.825 91.100 ;
        RECT 303.080 90.935 303.250 91.665 ;
        RECT 303.425 91.590 303.685 92.740 ;
        RECT 303.860 91.575 304.150 92.740 ;
        RECT 304.320 91.770 304.630 92.570 ;
        RECT 304.800 91.940 305.110 92.740 ;
        RECT 305.280 92.110 305.540 92.570 ;
        RECT 305.710 92.280 305.965 92.740 ;
        RECT 306.140 92.110 306.400 92.570 ;
        RECT 305.280 91.940 306.400 92.110 ;
        RECT 304.320 91.600 305.350 91.770 ;
        RECT 302.110 90.740 302.825 90.910 ;
        RECT 302.110 90.360 302.280 90.740 ;
        RECT 302.495 90.190 302.825 90.570 ;
        RECT 302.995 90.360 303.250 90.935 ;
        RECT 303.425 90.190 303.685 91.030 ;
        RECT 303.860 90.190 304.150 90.915 ;
        RECT 304.320 90.690 304.490 91.600 ;
        RECT 304.660 90.860 305.010 91.430 ;
        RECT 305.180 91.350 305.350 91.600 ;
        RECT 306.140 91.690 306.400 91.940 ;
        RECT 306.570 91.870 306.855 92.740 ;
        RECT 308.090 91.810 308.260 92.570 ;
        RECT 308.475 91.980 308.805 92.740 ;
        RECT 306.140 91.520 306.895 91.690 ;
        RECT 308.090 91.640 308.805 91.810 ;
        RECT 308.975 91.665 309.230 92.570 ;
        RECT 305.180 91.180 306.320 91.350 ;
        RECT 306.490 91.010 306.895 91.520 ;
        RECT 308.000 91.090 308.355 91.460 ;
        RECT 308.635 91.430 308.805 91.640 ;
        RECT 308.635 91.100 308.890 91.430 ;
        RECT 305.245 90.840 306.895 91.010 ;
        RECT 308.635 90.910 308.805 91.100 ;
        RECT 309.060 90.935 309.230 91.665 ;
        RECT 309.405 91.590 309.665 92.740 ;
        RECT 309.840 91.650 311.050 92.740 ;
        RECT 309.840 91.110 310.360 91.650 ;
        RECT 304.320 90.360 304.620 90.690 ;
        RECT 304.790 90.190 305.065 90.670 ;
        RECT 305.245 90.450 305.540 90.840 ;
        RECT 305.710 90.190 305.965 90.670 ;
        RECT 306.140 90.450 306.400 90.840 ;
        RECT 308.090 90.740 308.805 90.910 ;
        RECT 306.570 90.190 306.850 90.670 ;
        RECT 308.090 90.360 308.260 90.740 ;
        RECT 308.475 90.190 308.805 90.570 ;
        RECT 308.975 90.360 309.230 90.935 ;
        RECT 309.405 90.190 309.665 91.030 ;
        RECT 310.530 90.940 311.050 91.480 ;
        RECT 309.840 90.190 311.050 90.940 ;
        RECT 162.095 90.020 311.135 90.190 ;
        RECT 162.180 89.270 163.390 90.020 ;
        RECT 162.180 88.730 162.700 89.270 ;
        RECT 163.560 89.250 167.070 90.020 ;
        RECT 167.705 89.310 167.960 89.840 ;
        RECT 168.130 89.560 168.435 90.020 ;
        RECT 168.680 89.640 169.750 89.810 ;
        RECT 162.870 88.560 163.390 89.100 ;
        RECT 163.560 88.730 165.210 89.250 ;
        RECT 165.380 88.560 167.070 89.080 ;
        RECT 162.180 87.470 163.390 88.560 ;
        RECT 163.560 87.470 167.070 88.560 ;
        RECT 167.705 88.660 167.915 89.310 ;
        RECT 168.680 89.285 169.000 89.640 ;
        RECT 168.675 89.110 169.000 89.285 ;
        RECT 168.085 88.810 169.000 89.110 ;
        RECT 169.170 89.070 169.410 89.470 ;
        RECT 169.580 89.410 169.750 89.640 ;
        RECT 169.920 89.580 170.110 90.020 ;
        RECT 170.280 89.570 171.230 89.850 ;
        RECT 171.450 89.660 171.800 89.830 ;
        RECT 169.580 89.240 170.110 89.410 ;
        RECT 168.085 88.780 168.825 88.810 ;
        RECT 167.705 87.780 167.960 88.660 ;
        RECT 168.130 87.470 168.435 88.610 ;
        RECT 168.655 88.190 168.825 88.780 ;
        RECT 169.170 88.700 169.710 89.070 ;
        RECT 169.890 88.960 170.110 89.240 ;
        RECT 170.280 88.790 170.450 89.570 ;
        RECT 170.045 88.620 170.450 88.790 ;
        RECT 170.620 88.780 170.970 89.400 ;
        RECT 170.045 88.530 170.215 88.620 ;
        RECT 171.140 88.610 171.350 89.400 ;
        RECT 168.995 88.360 170.215 88.530 ;
        RECT 170.675 88.450 171.350 88.610 ;
        RECT 168.655 88.020 169.455 88.190 ;
        RECT 168.775 87.470 169.105 87.850 ;
        RECT 169.285 87.730 169.455 88.020 ;
        RECT 170.045 87.980 170.215 88.360 ;
        RECT 170.385 88.440 171.350 88.450 ;
        RECT 171.540 89.270 171.800 89.660 ;
        RECT 172.010 89.560 172.340 90.020 ;
        RECT 173.215 89.630 174.070 89.800 ;
        RECT 174.275 89.630 174.770 89.800 ;
        RECT 174.940 89.660 175.270 90.020 ;
        RECT 171.540 88.580 171.710 89.270 ;
        RECT 171.880 88.920 172.050 89.100 ;
        RECT 172.220 89.090 173.010 89.340 ;
        RECT 173.215 88.920 173.385 89.630 ;
        RECT 173.555 89.120 173.910 89.340 ;
        RECT 171.880 88.750 173.570 88.920 ;
        RECT 170.385 88.150 170.845 88.440 ;
        RECT 171.540 88.410 173.040 88.580 ;
        RECT 171.540 88.270 171.710 88.410 ;
        RECT 171.150 88.100 171.710 88.270 ;
        RECT 169.625 87.470 169.875 87.930 ;
        RECT 170.045 87.640 170.915 87.980 ;
        RECT 171.150 87.640 171.320 88.100 ;
        RECT 172.155 88.070 173.230 88.240 ;
        RECT 171.490 87.470 171.860 87.930 ;
        RECT 172.155 87.730 172.325 88.070 ;
        RECT 172.495 87.470 172.825 87.900 ;
        RECT 173.060 87.730 173.230 88.070 ;
        RECT 173.400 87.970 173.570 88.750 ;
        RECT 173.740 88.530 173.910 89.120 ;
        RECT 174.080 88.720 174.430 89.340 ;
        RECT 173.740 88.140 174.205 88.530 ;
        RECT 174.600 88.270 174.770 89.630 ;
        RECT 174.940 88.440 175.400 89.490 ;
        RECT 174.375 88.100 174.770 88.270 ;
        RECT 174.375 87.970 174.545 88.100 ;
        RECT 173.400 87.640 174.080 87.970 ;
        RECT 174.295 87.640 174.545 87.970 ;
        RECT 174.715 87.470 174.965 87.930 ;
        RECT 175.135 87.655 175.460 88.440 ;
        RECT 175.630 87.640 175.800 89.760 ;
        RECT 175.970 89.640 176.300 90.020 ;
        RECT 176.470 89.470 176.725 89.760 ;
        RECT 175.975 89.300 176.725 89.470 ;
        RECT 175.975 88.310 176.205 89.300 ;
        RECT 176.905 89.280 177.160 89.850 ;
        RECT 177.330 89.620 177.660 90.020 ;
        RECT 178.085 89.485 178.615 89.850 ;
        RECT 178.085 89.450 178.260 89.485 ;
        RECT 177.330 89.280 178.260 89.450 ;
        RECT 176.375 88.480 176.725 89.130 ;
        RECT 176.905 88.610 177.075 89.280 ;
        RECT 177.330 89.110 177.500 89.280 ;
        RECT 177.245 88.780 177.500 89.110 ;
        RECT 177.725 88.780 177.920 89.110 ;
        RECT 175.975 88.140 176.725 88.310 ;
        RECT 175.970 87.470 176.300 87.970 ;
        RECT 176.470 87.640 176.725 88.140 ;
        RECT 176.905 87.640 177.240 88.610 ;
        RECT 177.410 87.470 177.580 88.610 ;
        RECT 177.750 87.810 177.920 88.780 ;
        RECT 178.090 88.150 178.260 89.280 ;
        RECT 178.430 88.490 178.600 89.290 ;
        RECT 178.805 89.000 179.080 89.850 ;
        RECT 178.800 88.830 179.080 89.000 ;
        RECT 178.805 88.690 179.080 88.830 ;
        RECT 179.250 88.490 179.440 89.850 ;
        RECT 179.620 89.485 180.130 90.020 ;
        RECT 180.350 89.210 180.595 89.815 ;
        RECT 181.040 89.280 181.425 89.850 ;
        RECT 181.595 89.560 181.920 90.020 ;
        RECT 182.440 89.390 182.720 89.850 ;
        RECT 179.640 89.040 180.870 89.210 ;
        RECT 178.430 88.320 179.440 88.490 ;
        RECT 179.610 88.475 180.360 88.665 ;
        RECT 178.090 87.980 179.215 88.150 ;
        RECT 179.610 87.810 179.780 88.475 ;
        RECT 180.530 88.230 180.870 89.040 ;
        RECT 177.750 87.640 179.780 87.810 ;
        RECT 179.950 87.470 180.120 88.230 ;
        RECT 180.355 87.820 180.870 88.230 ;
        RECT 181.040 88.610 181.320 89.280 ;
        RECT 181.595 89.220 182.720 89.390 ;
        RECT 181.595 89.110 182.045 89.220 ;
        RECT 181.490 88.780 182.045 89.110 ;
        RECT 182.910 89.050 183.310 89.850 ;
        RECT 183.710 89.560 183.980 90.020 ;
        RECT 184.150 89.390 184.435 89.850 ;
        RECT 181.040 87.640 181.425 88.610 ;
        RECT 181.595 88.320 182.045 88.780 ;
        RECT 182.215 88.490 183.310 89.050 ;
        RECT 181.595 88.100 182.720 88.320 ;
        RECT 181.595 87.470 181.920 87.930 ;
        RECT 182.440 87.640 182.720 88.100 ;
        RECT 182.910 87.640 183.310 88.490 ;
        RECT 183.480 89.220 184.435 89.390 ;
        RECT 183.480 88.320 183.690 89.220 ;
        RECT 184.720 89.075 185.060 89.850 ;
        RECT 185.230 89.560 185.400 90.020 ;
        RECT 185.640 89.585 186.000 89.850 ;
        RECT 185.640 89.580 185.995 89.585 ;
        RECT 185.640 89.570 185.990 89.580 ;
        RECT 185.640 89.565 185.985 89.570 ;
        RECT 185.640 89.555 185.980 89.565 ;
        RECT 186.630 89.560 186.800 90.020 ;
        RECT 185.640 89.550 185.975 89.555 ;
        RECT 185.640 89.540 185.965 89.550 ;
        RECT 185.640 89.530 185.955 89.540 ;
        RECT 185.640 89.390 185.940 89.530 ;
        RECT 185.230 89.200 185.940 89.390 ;
        RECT 186.130 89.390 186.460 89.470 ;
        RECT 186.970 89.390 187.310 89.850 ;
        RECT 186.130 89.200 187.310 89.390 ;
        RECT 187.940 89.295 188.230 90.020 ;
        RECT 188.400 89.250 191.910 90.020 ;
        RECT 193.035 89.280 193.650 89.850 ;
        RECT 193.820 89.510 194.035 90.020 ;
        RECT 194.265 89.510 194.545 89.840 ;
        RECT 194.725 89.510 194.965 90.020 ;
        RECT 183.860 88.490 184.550 89.050 ;
        RECT 183.480 88.100 184.435 88.320 ;
        RECT 183.710 87.470 183.980 87.930 ;
        RECT 184.150 87.640 184.435 88.100 ;
        RECT 184.720 87.640 185.000 89.075 ;
        RECT 185.230 88.630 185.515 89.200 ;
        RECT 185.700 88.800 186.170 89.030 ;
        RECT 186.340 89.010 186.670 89.030 ;
        RECT 186.340 88.830 186.790 89.010 ;
        RECT 186.980 88.830 187.310 89.030 ;
        RECT 185.230 88.415 186.380 88.630 ;
        RECT 185.170 87.470 185.880 88.245 ;
        RECT 186.050 87.640 186.380 88.415 ;
        RECT 186.575 87.715 186.790 88.830 ;
        RECT 187.080 88.490 187.310 88.830 ;
        RECT 188.400 88.730 190.050 89.250 ;
        RECT 186.970 87.470 187.300 88.190 ;
        RECT 187.940 87.470 188.230 88.635 ;
        RECT 190.220 88.560 191.910 89.080 ;
        RECT 188.400 87.470 191.910 88.560 ;
        RECT 193.035 88.260 193.350 89.280 ;
        RECT 193.520 88.610 193.690 89.110 ;
        RECT 193.940 88.780 194.205 89.340 ;
        RECT 194.375 88.610 194.545 89.510 ;
        RECT 195.300 89.475 200.645 90.020 ;
        RECT 200.985 89.510 201.225 90.020 ;
        RECT 201.405 89.510 201.685 89.840 ;
        RECT 201.915 89.510 202.130 90.020 ;
        RECT 194.715 88.780 195.070 89.340 ;
        RECT 196.885 88.645 197.225 89.475 ;
        RECT 193.520 88.440 194.945 88.610 ;
        RECT 193.035 87.640 193.570 88.260 ;
        RECT 193.740 87.470 194.070 88.270 ;
        RECT 194.555 88.265 194.945 88.440 ;
        RECT 198.705 87.905 199.055 89.155 ;
        RECT 200.880 88.780 201.235 89.340 ;
        RECT 201.405 88.610 201.575 89.510 ;
        RECT 201.745 88.780 202.010 89.340 ;
        RECT 202.300 89.280 202.915 89.850 ;
        RECT 203.140 89.290 203.430 90.020 ;
        RECT 202.260 88.610 202.430 89.110 ;
        RECT 201.005 88.440 202.430 88.610 ;
        RECT 201.005 88.265 201.395 88.440 ;
        RECT 195.300 87.470 200.645 87.905 ;
        RECT 201.880 87.470 202.210 88.270 ;
        RECT 202.600 88.260 202.915 89.280 ;
        RECT 203.130 88.780 203.430 89.110 ;
        RECT 203.610 89.090 203.840 89.730 ;
        RECT 204.020 89.470 204.330 89.840 ;
        RECT 204.510 89.650 205.180 90.020 ;
        RECT 204.020 89.270 205.250 89.470 ;
        RECT 203.610 88.780 204.135 89.090 ;
        RECT 204.315 88.780 204.780 89.090 ;
        RECT 204.960 88.600 205.250 89.270 ;
        RECT 202.380 87.640 202.915 88.260 ;
        RECT 203.140 88.360 204.300 88.600 ;
        RECT 203.140 87.650 203.400 88.360 ;
        RECT 203.570 87.470 203.900 88.180 ;
        RECT 204.070 87.650 204.300 88.360 ;
        RECT 204.480 88.380 205.250 88.600 ;
        RECT 204.480 87.650 204.750 88.380 ;
        RECT 204.930 87.470 205.270 88.200 ;
        RECT 205.440 87.650 205.700 89.840 ;
        RECT 206.085 89.240 206.585 89.850 ;
        RECT 205.880 88.780 206.230 89.030 ;
        RECT 206.415 88.610 206.585 89.240 ;
        RECT 207.215 89.370 207.545 89.850 ;
        RECT 207.715 89.560 207.940 90.020 ;
        RECT 208.110 89.370 208.440 89.850 ;
        RECT 207.215 89.200 208.440 89.370 ;
        RECT 208.630 89.220 208.880 90.020 ;
        RECT 209.050 89.220 209.390 89.850 ;
        RECT 206.755 88.830 207.085 89.030 ;
        RECT 207.255 88.830 207.585 89.030 ;
        RECT 207.755 88.830 208.175 89.030 ;
        RECT 208.350 88.860 209.045 89.030 ;
        RECT 208.350 88.610 208.520 88.860 ;
        RECT 209.215 88.610 209.390 89.220 ;
        RECT 209.560 89.250 213.070 90.020 ;
        RECT 213.700 89.295 213.990 90.020 ;
        RECT 214.210 89.480 214.435 89.840 ;
        RECT 214.615 89.650 214.945 90.020 ;
        RECT 215.125 89.480 215.380 89.840 ;
        RECT 215.945 89.650 216.690 90.020 ;
        RECT 214.210 89.290 216.695 89.480 ;
        RECT 209.560 88.730 211.210 89.250 ;
        RECT 206.085 88.440 208.520 88.610 ;
        RECT 206.085 87.640 206.415 88.440 ;
        RECT 206.585 87.470 206.915 88.270 ;
        RECT 207.215 87.640 207.545 88.440 ;
        RECT 208.190 87.470 208.440 88.270 ;
        RECT 208.710 87.470 208.880 88.610 ;
        RECT 209.050 87.640 209.390 88.610 ;
        RECT 211.380 88.560 213.070 89.080 ;
        RECT 214.170 88.780 214.440 89.110 ;
        RECT 214.620 88.780 215.055 89.110 ;
        RECT 215.235 88.780 215.810 89.110 ;
        RECT 215.990 88.780 216.270 89.110 ;
        RECT 209.560 87.470 213.070 88.560 ;
        RECT 213.700 87.470 213.990 88.635 ;
        RECT 216.470 88.600 216.695 89.290 ;
        RECT 214.200 88.420 216.695 88.600 ;
        RECT 216.870 88.420 217.205 89.840 ;
        RECT 217.380 89.475 222.725 90.020 ;
        RECT 218.965 88.645 219.305 89.475 ;
        RECT 222.900 89.250 225.490 90.020 ;
        RECT 226.125 89.255 226.580 90.020 ;
        RECT 226.855 89.640 228.155 89.850 ;
        RECT 228.410 89.660 228.740 90.020 ;
        RECT 227.985 89.490 228.155 89.640 ;
        RECT 228.910 89.520 229.170 89.850 ;
        RECT 228.940 89.510 229.170 89.520 ;
        RECT 214.200 87.650 214.490 88.420 ;
        RECT 215.060 88.010 216.250 88.240 ;
        RECT 215.060 87.650 215.320 88.010 ;
        RECT 215.490 87.470 215.820 87.840 ;
        RECT 215.990 87.650 216.250 88.010 ;
        RECT 216.440 87.470 216.770 88.190 ;
        RECT 216.940 87.650 217.205 88.420 ;
        RECT 220.785 87.905 221.135 89.155 ;
        RECT 222.900 88.730 224.110 89.250 ;
        RECT 224.280 88.560 225.490 89.080 ;
        RECT 227.055 89.030 227.275 89.430 ;
        RECT 226.120 88.830 226.610 89.030 ;
        RECT 226.800 88.820 227.275 89.030 ;
        RECT 227.520 89.030 227.730 89.430 ;
        RECT 227.985 89.365 228.740 89.490 ;
        RECT 227.985 89.320 228.830 89.365 ;
        RECT 228.560 89.200 228.830 89.320 ;
        RECT 227.520 88.820 227.850 89.030 ;
        RECT 228.020 88.760 228.430 89.065 ;
        RECT 217.380 87.470 222.725 87.905 ;
        RECT 222.900 87.470 225.490 88.560 ;
        RECT 226.125 88.590 227.300 88.650 ;
        RECT 228.660 88.625 228.830 89.200 ;
        RECT 228.630 88.590 228.830 88.625 ;
        RECT 226.125 88.480 228.830 88.590 ;
        RECT 226.125 87.860 226.380 88.480 ;
        RECT 226.970 88.420 228.770 88.480 ;
        RECT 226.970 88.390 227.300 88.420 ;
        RECT 229.000 88.320 229.170 89.510 ;
        RECT 226.630 88.220 226.815 88.310 ;
        RECT 227.405 88.220 228.240 88.230 ;
        RECT 226.630 88.020 228.240 88.220 ;
        RECT 226.630 87.980 226.860 88.020 ;
        RECT 226.125 87.640 226.460 87.860 ;
        RECT 227.465 87.470 227.820 87.850 ;
        RECT 227.990 87.640 228.240 88.020 ;
        RECT 228.490 87.470 228.740 88.250 ;
        RECT 228.910 87.640 229.170 88.320 ;
        RECT 229.345 89.345 229.620 89.690 ;
        RECT 229.810 89.620 230.190 90.020 ;
        RECT 230.360 89.450 230.530 89.800 ;
        RECT 230.700 89.620 231.030 90.020 ;
        RECT 231.200 89.450 231.455 89.800 ;
        RECT 231.640 89.475 236.985 90.020 ;
        RECT 229.345 88.610 229.515 89.345 ;
        RECT 229.790 89.280 231.455 89.450 ;
        RECT 229.790 89.110 229.960 89.280 ;
        RECT 229.685 88.780 229.960 89.110 ;
        RECT 230.130 88.780 230.955 89.110 ;
        RECT 231.125 88.780 231.470 89.110 ;
        RECT 229.790 88.610 229.960 88.780 ;
        RECT 229.345 87.640 229.620 88.610 ;
        RECT 229.790 88.440 230.450 88.610 ;
        RECT 230.760 88.490 230.955 88.780 ;
        RECT 233.225 88.645 233.565 89.475 ;
        RECT 237.160 89.250 238.830 90.020 ;
        RECT 239.460 89.295 239.750 90.020 ;
        RECT 239.920 89.250 243.430 90.020 ;
        RECT 230.280 88.320 230.450 88.440 ;
        RECT 231.125 88.320 231.450 88.610 ;
        RECT 229.830 87.470 230.110 88.270 ;
        RECT 230.280 88.150 231.450 88.320 ;
        RECT 230.280 87.690 231.470 87.980 ;
        RECT 235.045 87.905 235.395 89.155 ;
        RECT 237.160 88.730 237.910 89.250 ;
        RECT 238.080 88.560 238.830 89.080 ;
        RECT 239.920 88.730 241.570 89.250 ;
        RECT 231.640 87.470 236.985 87.905 ;
        RECT 237.160 87.470 238.830 88.560 ;
        RECT 239.460 87.470 239.750 88.635 ;
        RECT 241.740 88.560 243.430 89.080 ;
        RECT 239.920 87.470 243.430 88.560 ;
        RECT 243.605 88.420 243.940 89.840 ;
        RECT 244.120 89.650 244.865 90.020 ;
        RECT 245.430 89.480 245.685 89.840 ;
        RECT 245.865 89.650 246.195 90.020 ;
        RECT 246.375 89.480 246.600 89.840 ;
        RECT 244.115 89.290 246.600 89.480 ;
        RECT 246.820 89.475 252.165 90.020 ;
        RECT 252.340 89.475 257.685 90.020 ;
        RECT 244.115 88.600 244.340 89.290 ;
        RECT 244.540 88.780 244.820 89.110 ;
        RECT 245.000 88.780 245.575 89.110 ;
        RECT 245.755 88.780 246.190 89.110 ;
        RECT 246.370 88.780 246.640 89.110 ;
        RECT 248.405 88.645 248.745 89.475 ;
        RECT 244.115 88.420 246.610 88.600 ;
        RECT 243.605 87.650 243.870 88.420 ;
        RECT 244.040 87.470 244.370 88.190 ;
        RECT 244.560 88.010 245.750 88.240 ;
        RECT 244.560 87.650 244.820 88.010 ;
        RECT 244.990 87.470 245.320 87.840 ;
        RECT 245.490 87.650 245.750 88.010 ;
        RECT 246.320 87.650 246.610 88.420 ;
        RECT 250.225 87.905 250.575 89.155 ;
        RECT 253.925 88.645 254.265 89.475 ;
        RECT 257.860 89.250 260.450 90.020 ;
        RECT 261.170 89.370 261.340 89.850 ;
        RECT 261.510 89.540 261.840 90.020 ;
        RECT 262.065 89.600 263.600 89.850 ;
        RECT 262.065 89.370 262.235 89.600 ;
        RECT 255.745 87.905 256.095 89.155 ;
        RECT 257.860 88.730 259.070 89.250 ;
        RECT 261.170 89.200 262.235 89.370 ;
        RECT 259.240 88.560 260.450 89.080 ;
        RECT 262.415 89.030 262.695 89.430 ;
        RECT 261.085 88.820 261.435 89.030 ;
        RECT 261.605 88.830 262.050 89.030 ;
        RECT 262.220 88.830 262.695 89.030 ;
        RECT 262.965 89.030 263.250 89.430 ;
        RECT 263.430 89.370 263.600 89.600 ;
        RECT 263.770 89.540 264.100 90.020 ;
        RECT 264.315 89.520 264.570 89.850 ;
        RECT 264.385 89.440 264.570 89.520 ;
        RECT 263.430 89.200 264.230 89.370 ;
        RECT 262.965 88.830 263.295 89.030 ;
        RECT 263.465 89.000 263.830 89.030 ;
        RECT 263.465 88.830 263.840 89.000 ;
        RECT 264.060 88.650 264.230 89.200 ;
        RECT 246.820 87.470 252.165 87.905 ;
        RECT 252.340 87.470 257.685 87.905 ;
        RECT 257.860 87.470 260.450 88.560 ;
        RECT 261.170 88.480 264.230 88.650 ;
        RECT 261.170 87.640 261.340 88.480 ;
        RECT 264.400 88.320 264.570 89.440 ;
        RECT 265.220 89.295 265.510 90.020 ;
        RECT 265.685 89.255 266.140 90.020 ;
        RECT 266.415 89.640 267.715 89.850 ;
        RECT 267.970 89.660 268.300 90.020 ;
        RECT 267.545 89.490 267.715 89.640 ;
        RECT 268.470 89.520 268.730 89.850 ;
        RECT 268.500 89.510 268.730 89.520 ;
        RECT 266.615 89.030 266.835 89.430 ;
        RECT 265.680 88.830 266.170 89.030 ;
        RECT 266.360 88.820 266.835 89.030 ;
        RECT 267.080 89.030 267.290 89.430 ;
        RECT 267.545 89.365 268.300 89.490 ;
        RECT 267.545 89.320 268.390 89.365 ;
        RECT 268.120 89.200 268.390 89.320 ;
        RECT 267.080 88.820 267.410 89.030 ;
        RECT 267.580 88.760 267.990 89.065 ;
        RECT 264.360 88.310 264.570 88.320 ;
        RECT 261.510 87.810 261.840 88.310 ;
        RECT 262.010 88.070 263.645 88.310 ;
        RECT 262.010 87.980 262.240 88.070 ;
        RECT 262.350 87.810 262.680 87.850 ;
        RECT 261.510 87.640 262.680 87.810 ;
        RECT 262.870 87.470 263.225 87.890 ;
        RECT 263.395 87.640 263.645 88.070 ;
        RECT 263.815 87.470 264.145 88.230 ;
        RECT 264.315 87.640 264.570 88.310 ;
        RECT 265.220 87.470 265.510 88.635 ;
        RECT 265.685 88.590 266.860 88.650 ;
        RECT 268.220 88.625 268.390 89.200 ;
        RECT 268.190 88.590 268.390 88.625 ;
        RECT 265.685 88.480 268.390 88.590 ;
        RECT 265.685 87.860 265.940 88.480 ;
        RECT 266.530 88.420 268.330 88.480 ;
        RECT 266.530 88.390 266.860 88.420 ;
        RECT 268.560 88.320 268.730 89.510 ;
        RECT 268.915 89.450 269.170 89.800 ;
        RECT 269.340 89.620 269.670 90.020 ;
        RECT 269.840 89.450 270.010 89.800 ;
        RECT 270.180 89.620 270.560 90.020 ;
        RECT 268.915 89.280 270.580 89.450 ;
        RECT 270.750 89.345 271.025 89.690 ;
        RECT 271.200 89.475 276.545 90.020 ;
        RECT 270.410 89.110 270.580 89.280 ;
        RECT 268.900 88.780 269.245 89.110 ;
        RECT 269.415 88.780 270.240 89.110 ;
        RECT 270.410 88.780 270.685 89.110 ;
        RECT 266.190 88.220 266.375 88.310 ;
        RECT 266.965 88.220 267.800 88.230 ;
        RECT 266.190 88.020 267.800 88.220 ;
        RECT 266.190 87.980 266.420 88.020 ;
        RECT 265.685 87.640 266.020 87.860 ;
        RECT 267.025 87.470 267.380 87.850 ;
        RECT 267.550 87.640 267.800 88.020 ;
        RECT 268.050 87.470 268.300 88.250 ;
        RECT 268.470 87.640 268.730 88.320 ;
        RECT 268.920 88.320 269.245 88.610 ;
        RECT 269.415 88.490 269.610 88.780 ;
        RECT 270.410 88.610 270.580 88.780 ;
        RECT 270.855 88.610 271.025 89.345 ;
        RECT 272.785 88.645 273.125 89.475 ;
        RECT 276.720 89.270 277.930 90.020 ;
        RECT 278.110 89.520 278.440 90.020 ;
        RECT 278.640 89.450 278.810 89.800 ;
        RECT 279.010 89.620 279.340 90.020 ;
        RECT 279.510 89.450 279.680 89.800 ;
        RECT 279.850 89.620 280.230 90.020 ;
        RECT 269.920 88.440 270.580 88.610 ;
        RECT 269.920 88.320 270.090 88.440 ;
        RECT 268.920 88.150 270.090 88.320 ;
        RECT 268.900 87.690 270.090 87.980 ;
        RECT 270.260 87.470 270.540 88.270 ;
        RECT 270.750 87.640 271.025 88.610 ;
        RECT 274.605 87.905 274.955 89.155 ;
        RECT 276.720 88.730 277.240 89.270 ;
        RECT 277.410 88.560 277.930 89.100 ;
        RECT 278.105 88.780 278.455 89.350 ;
        RECT 278.640 89.280 280.250 89.450 ;
        RECT 280.420 89.345 280.690 89.690 ;
        RECT 280.860 89.475 286.205 90.020 ;
        RECT 280.080 89.110 280.250 89.280 ;
        RECT 271.200 87.470 276.545 87.905 ;
        RECT 276.720 87.470 277.930 88.560 ;
        RECT 278.105 88.320 278.425 88.610 ;
        RECT 278.625 88.490 279.335 89.110 ;
        RECT 279.505 88.780 279.910 89.110 ;
        RECT 280.080 88.780 280.350 89.110 ;
        RECT 280.080 88.610 280.250 88.780 ;
        RECT 280.520 88.610 280.690 89.345 ;
        RECT 282.445 88.645 282.785 89.475 ;
        RECT 286.380 89.250 289.890 90.020 ;
        RECT 290.980 89.295 291.270 90.020 ;
        RECT 291.440 89.250 294.950 90.020 ;
        RECT 295.125 89.470 295.380 89.760 ;
        RECT 295.550 89.640 295.880 90.020 ;
        RECT 295.125 89.300 295.875 89.470 ;
        RECT 279.525 88.440 280.250 88.610 ;
        RECT 279.525 88.320 279.695 88.440 ;
        RECT 278.105 88.150 279.695 88.320 ;
        RECT 278.105 87.690 279.760 87.980 ;
        RECT 279.930 87.470 280.210 88.270 ;
        RECT 280.420 87.640 280.690 88.610 ;
        RECT 284.265 87.905 284.615 89.155 ;
        RECT 286.380 88.730 288.030 89.250 ;
        RECT 288.200 88.560 289.890 89.080 ;
        RECT 291.440 88.730 293.090 89.250 ;
        RECT 280.860 87.470 286.205 87.905 ;
        RECT 286.380 87.470 289.890 88.560 ;
        RECT 290.980 87.470 291.270 88.635 ;
        RECT 293.260 88.560 294.950 89.080 ;
        RECT 291.440 87.470 294.950 88.560 ;
        RECT 295.125 88.480 295.475 89.130 ;
        RECT 295.645 88.310 295.875 89.300 ;
        RECT 295.125 88.140 295.875 88.310 ;
        RECT 295.125 87.640 295.380 88.140 ;
        RECT 295.550 87.470 295.880 87.970 ;
        RECT 296.050 87.640 296.220 89.760 ;
        RECT 296.580 89.660 296.910 90.020 ;
        RECT 297.080 89.630 297.575 89.800 ;
        RECT 297.780 89.630 298.635 89.800 ;
        RECT 296.450 88.440 296.910 89.490 ;
        RECT 296.390 87.655 296.715 88.440 ;
        RECT 297.080 88.270 297.250 89.630 ;
        RECT 297.420 88.720 297.770 89.340 ;
        RECT 297.940 89.120 298.295 89.340 ;
        RECT 297.940 88.530 298.110 89.120 ;
        RECT 298.465 88.920 298.635 89.630 ;
        RECT 299.510 89.560 299.840 90.020 ;
        RECT 300.050 89.660 300.400 89.830 ;
        RECT 298.840 89.090 299.630 89.340 ;
        RECT 300.050 89.270 300.310 89.660 ;
        RECT 300.620 89.570 301.570 89.850 ;
        RECT 301.740 89.580 301.930 90.020 ;
        RECT 302.100 89.640 303.170 89.810 ;
        RECT 299.800 88.920 299.970 89.100 ;
        RECT 297.080 88.100 297.475 88.270 ;
        RECT 297.645 88.140 298.110 88.530 ;
        RECT 298.280 88.750 299.970 88.920 ;
        RECT 297.305 87.970 297.475 88.100 ;
        RECT 298.280 87.970 298.450 88.750 ;
        RECT 300.140 88.580 300.310 89.270 ;
        RECT 298.810 88.410 300.310 88.580 ;
        RECT 300.500 88.610 300.710 89.400 ;
        RECT 300.880 88.780 301.230 89.400 ;
        RECT 301.400 88.790 301.570 89.570 ;
        RECT 302.100 89.410 302.270 89.640 ;
        RECT 301.740 89.240 302.270 89.410 ;
        RECT 301.740 88.960 301.960 89.240 ;
        RECT 302.440 89.070 302.680 89.470 ;
        RECT 301.400 88.620 301.805 88.790 ;
        RECT 302.140 88.700 302.680 89.070 ;
        RECT 302.850 89.285 303.170 89.640 ;
        RECT 303.415 89.560 303.720 90.020 ;
        RECT 303.890 89.310 304.140 89.840 ;
        RECT 302.850 89.110 303.175 89.285 ;
        RECT 302.850 88.810 303.765 89.110 ;
        RECT 303.025 88.780 303.765 88.810 ;
        RECT 300.500 88.450 301.175 88.610 ;
        RECT 301.635 88.530 301.805 88.620 ;
        RECT 300.500 88.440 301.465 88.450 ;
        RECT 300.140 88.270 300.310 88.410 ;
        RECT 296.885 87.470 297.135 87.930 ;
        RECT 297.305 87.640 297.555 87.970 ;
        RECT 297.770 87.640 298.450 87.970 ;
        RECT 298.620 88.070 299.695 88.240 ;
        RECT 300.140 88.100 300.700 88.270 ;
        RECT 301.005 88.150 301.465 88.440 ;
        RECT 301.635 88.360 302.855 88.530 ;
        RECT 298.620 87.730 298.790 88.070 ;
        RECT 299.025 87.470 299.355 87.900 ;
        RECT 299.525 87.730 299.695 88.070 ;
        RECT 299.990 87.470 300.360 87.930 ;
        RECT 300.530 87.640 300.700 88.100 ;
        RECT 301.635 87.980 301.805 88.360 ;
        RECT 303.025 88.190 303.195 88.780 ;
        RECT 303.935 88.660 304.140 89.310 ;
        RECT 304.310 89.265 304.560 90.020 ;
        RECT 304.780 89.270 305.990 90.020 ;
        RECT 306.250 89.470 306.420 89.850 ;
        RECT 306.635 89.640 306.965 90.020 ;
        RECT 306.250 89.300 306.965 89.470 ;
        RECT 304.780 88.730 305.300 89.270 ;
        RECT 300.935 87.640 301.805 87.980 ;
        RECT 302.395 88.020 303.195 88.190 ;
        RECT 301.975 87.470 302.225 87.930 ;
        RECT 302.395 87.730 302.565 88.020 ;
        RECT 302.745 87.470 303.075 87.850 ;
        RECT 303.415 87.470 303.720 88.610 ;
        RECT 303.890 87.780 304.140 88.660 ;
        RECT 304.310 87.470 304.560 88.610 ;
        RECT 305.470 88.560 305.990 89.100 ;
        RECT 306.160 88.750 306.515 89.120 ;
        RECT 306.795 89.110 306.965 89.300 ;
        RECT 307.135 89.275 307.390 89.850 ;
        RECT 306.795 88.780 307.050 89.110 ;
        RECT 306.795 88.570 306.965 88.780 ;
        RECT 304.780 87.470 305.990 88.560 ;
        RECT 306.250 88.400 306.965 88.570 ;
        RECT 307.220 88.545 307.390 89.275 ;
        RECT 307.565 89.180 307.825 90.020 ;
        RECT 308.090 89.470 308.260 89.850 ;
        RECT 308.475 89.640 308.805 90.020 ;
        RECT 308.090 89.300 308.805 89.470 ;
        RECT 308.000 88.750 308.355 89.120 ;
        RECT 308.635 89.110 308.805 89.300 ;
        RECT 308.975 89.275 309.230 89.850 ;
        RECT 308.635 88.780 308.890 89.110 ;
        RECT 306.250 87.640 306.420 88.400 ;
        RECT 306.635 87.470 306.965 88.230 ;
        RECT 307.135 87.640 307.390 88.545 ;
        RECT 307.565 87.470 307.825 88.620 ;
        RECT 308.635 88.570 308.805 88.780 ;
        RECT 308.090 88.400 308.805 88.570 ;
        RECT 309.060 88.545 309.230 89.275 ;
        RECT 309.405 89.180 309.665 90.020 ;
        RECT 309.840 89.270 311.050 90.020 ;
        RECT 308.090 87.640 308.260 88.400 ;
        RECT 308.475 87.470 308.805 88.230 ;
        RECT 308.975 87.640 309.230 88.545 ;
        RECT 309.405 87.470 309.665 88.620 ;
        RECT 309.840 88.560 310.360 89.100 ;
        RECT 310.530 88.730 311.050 89.270 ;
        RECT 309.840 87.470 311.050 88.560 ;
        RECT 162.095 87.300 311.135 87.470 ;
        RECT 162.180 86.210 163.390 87.300 ;
        RECT 163.560 86.210 165.230 87.300 ;
        RECT 165.865 86.630 166.120 87.130 ;
        RECT 166.290 86.800 166.620 87.300 ;
        RECT 165.865 86.460 166.615 86.630 ;
        RECT 162.180 85.500 162.700 86.040 ;
        RECT 162.870 85.670 163.390 86.210 ;
        RECT 163.560 85.520 164.310 86.040 ;
        RECT 164.480 85.690 165.230 86.210 ;
        RECT 165.865 85.640 166.215 86.290 ;
        RECT 162.180 84.750 163.390 85.500 ;
        RECT 163.560 84.750 165.230 85.520 ;
        RECT 166.385 85.470 166.615 86.460 ;
        RECT 165.865 85.300 166.615 85.470 ;
        RECT 165.865 85.010 166.120 85.300 ;
        RECT 166.290 84.750 166.620 85.130 ;
        RECT 166.790 85.010 166.960 87.130 ;
        RECT 167.130 86.330 167.455 87.115 ;
        RECT 167.625 86.840 167.875 87.300 ;
        RECT 168.045 86.800 168.295 87.130 ;
        RECT 168.510 86.800 169.190 87.130 ;
        RECT 168.045 86.670 168.215 86.800 ;
        RECT 167.820 86.500 168.215 86.670 ;
        RECT 167.190 85.280 167.650 86.330 ;
        RECT 167.820 85.140 167.990 86.500 ;
        RECT 168.385 86.240 168.850 86.630 ;
        RECT 168.160 85.430 168.510 86.050 ;
        RECT 168.680 85.650 168.850 86.240 ;
        RECT 169.020 86.020 169.190 86.800 ;
        RECT 169.360 86.700 169.530 87.040 ;
        RECT 169.765 86.870 170.095 87.300 ;
        RECT 170.265 86.700 170.435 87.040 ;
        RECT 170.730 86.840 171.100 87.300 ;
        RECT 169.360 86.530 170.435 86.700 ;
        RECT 171.270 86.670 171.440 87.130 ;
        RECT 171.675 86.790 172.545 87.130 ;
        RECT 172.715 86.840 172.965 87.300 ;
        RECT 170.880 86.500 171.440 86.670 ;
        RECT 170.880 86.360 171.050 86.500 ;
        RECT 169.550 86.190 171.050 86.360 ;
        RECT 171.745 86.330 172.205 86.620 ;
        RECT 169.020 85.850 170.710 86.020 ;
        RECT 168.680 85.430 169.035 85.650 ;
        RECT 169.205 85.140 169.375 85.850 ;
        RECT 169.580 85.430 170.370 85.680 ;
        RECT 170.540 85.670 170.710 85.850 ;
        RECT 170.880 85.500 171.050 86.190 ;
        RECT 167.320 84.750 167.650 85.110 ;
        RECT 167.820 84.970 168.315 85.140 ;
        RECT 168.520 84.970 169.375 85.140 ;
        RECT 170.250 84.750 170.580 85.210 ;
        RECT 170.790 85.110 171.050 85.500 ;
        RECT 171.240 86.320 172.205 86.330 ;
        RECT 172.375 86.410 172.545 86.790 ;
        RECT 173.135 86.750 173.305 87.040 ;
        RECT 173.485 86.920 173.815 87.300 ;
        RECT 173.135 86.580 173.935 86.750 ;
        RECT 171.240 86.160 171.915 86.320 ;
        RECT 172.375 86.240 173.595 86.410 ;
        RECT 171.240 85.370 171.450 86.160 ;
        RECT 172.375 86.150 172.545 86.240 ;
        RECT 171.620 85.370 171.970 85.990 ;
        RECT 172.140 85.980 172.545 86.150 ;
        RECT 172.140 85.200 172.310 85.980 ;
        RECT 172.480 85.530 172.700 85.810 ;
        RECT 172.880 85.700 173.420 86.070 ;
        RECT 173.765 85.990 173.935 86.580 ;
        RECT 174.155 86.160 174.460 87.300 ;
        RECT 174.630 86.110 174.885 86.990 ;
        RECT 175.060 86.135 175.350 87.300 ;
        RECT 175.525 86.630 175.780 87.130 ;
        RECT 175.950 86.800 176.280 87.300 ;
        RECT 175.525 86.460 176.275 86.630 ;
        RECT 173.765 85.960 174.505 85.990 ;
        RECT 172.480 85.360 173.010 85.530 ;
        RECT 170.790 84.940 171.140 85.110 ;
        RECT 171.360 84.920 172.310 85.200 ;
        RECT 172.480 84.750 172.670 85.190 ;
        RECT 172.840 85.130 173.010 85.360 ;
        RECT 173.180 85.300 173.420 85.700 ;
        RECT 173.590 85.660 174.505 85.960 ;
        RECT 173.590 85.485 173.915 85.660 ;
        RECT 173.590 85.130 173.910 85.485 ;
        RECT 174.675 85.460 174.885 86.110 ;
        RECT 175.525 85.640 175.875 86.290 ;
        RECT 172.840 84.960 173.910 85.130 ;
        RECT 174.155 84.750 174.460 85.210 ;
        RECT 174.630 84.930 174.885 85.460 ;
        RECT 175.060 84.750 175.350 85.475 ;
        RECT 176.045 85.470 176.275 86.460 ;
        RECT 175.525 85.300 176.275 85.470 ;
        RECT 175.525 85.010 175.780 85.300 ;
        RECT 175.950 84.750 176.280 85.130 ;
        RECT 176.450 85.010 176.620 87.130 ;
        RECT 176.790 86.330 177.115 87.115 ;
        RECT 177.285 86.840 177.535 87.300 ;
        RECT 177.705 86.800 177.955 87.130 ;
        RECT 178.170 86.800 178.850 87.130 ;
        RECT 177.705 86.670 177.875 86.800 ;
        RECT 177.480 86.500 177.875 86.670 ;
        RECT 176.850 85.280 177.310 86.330 ;
        RECT 177.480 85.140 177.650 86.500 ;
        RECT 178.045 86.240 178.510 86.630 ;
        RECT 177.820 85.430 178.170 86.050 ;
        RECT 178.340 85.650 178.510 86.240 ;
        RECT 178.680 86.020 178.850 86.800 ;
        RECT 179.020 86.700 179.190 87.040 ;
        RECT 179.425 86.870 179.755 87.300 ;
        RECT 179.925 86.700 180.095 87.040 ;
        RECT 180.390 86.840 180.760 87.300 ;
        RECT 179.020 86.530 180.095 86.700 ;
        RECT 180.930 86.670 181.100 87.130 ;
        RECT 181.335 86.790 182.205 87.130 ;
        RECT 182.375 86.840 182.625 87.300 ;
        RECT 180.540 86.500 181.100 86.670 ;
        RECT 180.540 86.360 180.710 86.500 ;
        RECT 179.210 86.190 180.710 86.360 ;
        RECT 181.405 86.330 181.865 86.620 ;
        RECT 178.680 85.850 180.370 86.020 ;
        RECT 178.340 85.430 178.695 85.650 ;
        RECT 178.865 85.140 179.035 85.850 ;
        RECT 179.240 85.430 180.030 85.680 ;
        RECT 180.200 85.670 180.370 85.850 ;
        RECT 180.540 85.500 180.710 86.190 ;
        RECT 176.980 84.750 177.310 85.110 ;
        RECT 177.480 84.970 177.975 85.140 ;
        RECT 178.180 84.970 179.035 85.140 ;
        RECT 179.910 84.750 180.240 85.210 ;
        RECT 180.450 85.110 180.710 85.500 ;
        RECT 180.900 86.320 181.865 86.330 ;
        RECT 182.035 86.410 182.205 86.790 ;
        RECT 182.795 86.750 182.965 87.040 ;
        RECT 183.145 86.920 183.475 87.300 ;
        RECT 182.795 86.580 183.595 86.750 ;
        RECT 180.900 86.160 181.575 86.320 ;
        RECT 182.035 86.240 183.255 86.410 ;
        RECT 180.900 85.370 181.110 86.160 ;
        RECT 182.035 86.150 182.205 86.240 ;
        RECT 181.280 85.370 181.630 85.990 ;
        RECT 181.800 85.980 182.205 86.150 ;
        RECT 181.800 85.200 181.970 85.980 ;
        RECT 182.140 85.530 182.360 85.810 ;
        RECT 182.540 85.700 183.080 86.070 ;
        RECT 183.425 85.990 183.595 86.580 ;
        RECT 183.815 86.160 184.120 87.300 ;
        RECT 184.290 86.110 184.545 86.990 ;
        RECT 184.720 86.160 185.010 87.300 ;
        RECT 185.180 86.580 185.630 87.130 ;
        RECT 185.820 86.580 186.150 87.300 ;
        RECT 183.425 85.960 184.165 85.990 ;
        RECT 182.140 85.360 182.670 85.530 ;
        RECT 180.450 84.940 180.800 85.110 ;
        RECT 181.020 84.920 181.970 85.200 ;
        RECT 182.140 84.750 182.330 85.190 ;
        RECT 182.500 85.130 182.670 85.360 ;
        RECT 182.840 85.300 183.080 85.700 ;
        RECT 183.250 85.660 184.165 85.960 ;
        RECT 183.250 85.485 183.575 85.660 ;
        RECT 183.250 85.130 183.570 85.485 ;
        RECT 184.335 85.460 184.545 86.110 ;
        RECT 182.500 84.960 183.570 85.130 ;
        RECT 183.815 84.750 184.120 85.210 ;
        RECT 184.290 84.930 184.545 85.460 ;
        RECT 184.720 84.750 185.010 85.550 ;
        RECT 185.180 85.210 185.430 86.580 ;
        RECT 186.360 86.410 186.660 86.960 ;
        RECT 186.830 86.630 187.110 87.300 ;
        RECT 185.720 86.240 186.660 86.410 ;
        RECT 185.720 85.990 185.890 86.240 ;
        RECT 186.995 85.990 187.310 86.430 ;
        RECT 187.480 86.160 187.770 87.300 ;
        RECT 187.940 86.580 188.390 87.130 ;
        RECT 188.580 86.580 188.910 87.300 ;
        RECT 185.600 85.660 185.890 85.990 ;
        RECT 186.060 85.740 186.390 85.990 ;
        RECT 186.620 85.740 187.310 85.990 ;
        RECT 185.720 85.570 185.890 85.660 ;
        RECT 185.720 85.380 187.110 85.570 ;
        RECT 185.180 84.920 185.730 85.210 ;
        RECT 185.900 84.750 186.150 85.210 ;
        RECT 186.780 85.020 187.110 85.380 ;
        RECT 187.480 84.750 187.770 85.550 ;
        RECT 187.940 85.210 188.190 86.580 ;
        RECT 189.120 86.410 189.420 86.960 ;
        RECT 189.590 86.630 189.870 87.300 ;
        RECT 188.480 86.240 189.420 86.410 ;
        RECT 188.480 85.990 188.650 86.240 ;
        RECT 189.755 85.990 190.070 86.430 ;
        RECT 190.240 86.210 191.910 87.300 ;
        RECT 188.360 85.660 188.650 85.990 ;
        RECT 188.820 85.740 189.150 85.990 ;
        RECT 189.380 85.740 190.070 85.990 ;
        RECT 188.480 85.570 188.650 85.660 ;
        RECT 188.480 85.380 189.870 85.570 ;
        RECT 187.940 84.920 188.490 85.210 ;
        RECT 188.660 84.750 188.910 85.210 ;
        RECT 189.540 85.020 189.870 85.380 ;
        RECT 190.240 85.520 190.990 86.040 ;
        RECT 191.160 85.690 191.910 86.210 ;
        RECT 192.575 86.510 193.110 87.130 ;
        RECT 190.240 84.750 191.910 85.520 ;
        RECT 192.575 85.490 192.890 86.510 ;
        RECT 193.280 86.500 193.610 87.300 ;
        RECT 194.095 86.330 194.485 86.505 ;
        RECT 193.060 86.160 194.485 86.330 ;
        RECT 195.045 86.330 195.375 87.130 ;
        RECT 195.545 86.500 195.875 87.300 ;
        RECT 196.175 86.330 196.505 87.130 ;
        RECT 197.150 86.500 197.400 87.300 ;
        RECT 195.045 86.160 197.480 86.330 ;
        RECT 197.670 86.160 197.840 87.300 ;
        RECT 198.010 86.160 198.350 87.130 ;
        RECT 198.520 86.210 200.190 87.300 ;
        RECT 193.060 85.660 193.230 86.160 ;
        RECT 192.575 84.920 193.190 85.490 ;
        RECT 193.480 85.430 193.745 85.990 ;
        RECT 193.915 85.260 194.085 86.160 ;
        RECT 194.255 85.430 194.610 85.990 ;
        RECT 194.840 85.740 195.190 85.990 ;
        RECT 195.375 85.530 195.545 86.160 ;
        RECT 195.715 85.740 196.045 85.940 ;
        RECT 196.215 85.740 196.545 85.940 ;
        RECT 196.715 85.740 197.135 85.940 ;
        RECT 197.310 85.910 197.480 86.160 ;
        RECT 197.310 85.740 198.005 85.910 ;
        RECT 193.360 84.750 193.575 85.260 ;
        RECT 193.805 84.930 194.085 85.260 ;
        RECT 194.265 84.750 194.505 85.260 ;
        RECT 195.045 84.920 195.545 85.530 ;
        RECT 196.175 85.400 197.400 85.570 ;
        RECT 198.175 85.550 198.350 86.160 ;
        RECT 196.175 84.920 196.505 85.400 ;
        RECT 196.675 84.750 196.900 85.210 ;
        RECT 197.070 84.920 197.400 85.400 ;
        RECT 197.590 84.750 197.840 85.550 ;
        RECT 198.010 84.920 198.350 85.550 ;
        RECT 198.520 85.520 199.270 86.040 ;
        RECT 199.440 85.690 200.190 86.210 ;
        RECT 200.820 86.135 201.110 87.300 ;
        RECT 201.465 86.330 201.855 86.505 ;
        RECT 202.340 86.500 202.670 87.300 ;
        RECT 202.840 86.510 203.375 87.130 ;
        RECT 201.465 86.160 202.890 86.330 ;
        RECT 198.520 84.750 200.190 85.520 ;
        RECT 200.820 84.750 201.110 85.475 ;
        RECT 201.340 85.430 201.695 85.990 ;
        RECT 201.865 85.260 202.035 86.160 ;
        RECT 202.205 85.430 202.470 85.990 ;
        RECT 202.720 85.660 202.890 86.160 ;
        RECT 203.060 85.490 203.375 86.510 ;
        RECT 204.245 86.330 204.575 87.130 ;
        RECT 204.745 86.500 205.075 87.300 ;
        RECT 205.375 86.330 205.705 87.130 ;
        RECT 206.350 86.500 206.600 87.300 ;
        RECT 204.245 86.160 206.680 86.330 ;
        RECT 206.870 86.160 207.040 87.300 ;
        RECT 207.210 86.160 207.550 87.130 ;
        RECT 208.365 86.330 208.755 86.505 ;
        RECT 209.240 86.500 209.570 87.300 ;
        RECT 209.740 86.510 210.275 87.130 ;
        RECT 208.365 86.160 209.790 86.330 ;
        RECT 204.040 85.740 204.390 85.990 ;
        RECT 204.575 85.530 204.745 86.160 ;
        RECT 204.915 85.740 205.245 85.940 ;
        RECT 205.415 85.740 205.745 85.940 ;
        RECT 205.915 85.740 206.335 85.940 ;
        RECT 206.510 85.910 206.680 86.160 ;
        RECT 206.510 85.740 207.205 85.910 ;
        RECT 201.445 84.750 201.685 85.260 ;
        RECT 201.865 84.930 202.145 85.260 ;
        RECT 202.375 84.750 202.590 85.260 ;
        RECT 202.760 84.920 203.375 85.490 ;
        RECT 204.245 84.920 204.745 85.530 ;
        RECT 205.375 85.400 206.600 85.570 ;
        RECT 207.375 85.550 207.550 86.160 ;
        RECT 205.375 84.920 205.705 85.400 ;
        RECT 205.875 84.750 206.100 85.210 ;
        RECT 206.270 84.920 206.600 85.400 ;
        RECT 206.790 84.750 207.040 85.550 ;
        RECT 207.210 84.920 207.550 85.550 ;
        RECT 208.240 85.430 208.595 85.990 ;
        RECT 208.765 85.260 208.935 86.160 ;
        RECT 209.105 85.430 209.370 85.990 ;
        RECT 209.620 85.660 209.790 86.160 ;
        RECT 209.960 85.490 210.275 86.510 ;
        RECT 210.685 86.330 211.015 87.130 ;
        RECT 211.185 86.500 211.515 87.300 ;
        RECT 211.815 86.330 212.145 87.130 ;
        RECT 212.790 86.500 213.040 87.300 ;
        RECT 210.685 86.160 213.120 86.330 ;
        RECT 213.310 86.160 213.480 87.300 ;
        RECT 213.650 86.160 213.990 87.130 ;
        RECT 214.160 86.865 219.505 87.300 ;
        RECT 219.680 86.865 225.025 87.300 ;
        RECT 210.480 85.740 210.830 85.990 ;
        RECT 211.015 85.530 211.185 86.160 ;
        RECT 211.355 85.740 211.685 85.940 ;
        RECT 211.855 85.740 212.185 85.940 ;
        RECT 212.355 85.740 212.775 85.940 ;
        RECT 212.950 85.910 213.120 86.160 ;
        RECT 212.950 85.740 213.645 85.910 ;
        RECT 208.345 84.750 208.585 85.260 ;
        RECT 208.765 84.930 209.045 85.260 ;
        RECT 209.275 84.750 209.490 85.260 ;
        RECT 209.660 84.920 210.275 85.490 ;
        RECT 210.685 84.920 211.185 85.530 ;
        RECT 211.815 85.400 213.040 85.570 ;
        RECT 213.815 85.550 213.990 86.160 ;
        RECT 211.815 84.920 212.145 85.400 ;
        RECT 212.315 84.750 212.540 85.210 ;
        RECT 212.710 84.920 213.040 85.400 ;
        RECT 213.230 84.750 213.480 85.550 ;
        RECT 213.650 84.920 213.990 85.550 ;
        RECT 215.745 85.295 216.085 86.125 ;
        RECT 217.565 85.615 217.915 86.865 ;
        RECT 221.265 85.295 221.605 86.125 ;
        RECT 223.085 85.615 223.435 86.865 ;
        RECT 225.200 86.210 226.410 87.300 ;
        RECT 225.200 85.500 225.720 86.040 ;
        RECT 225.890 85.670 226.410 86.210 ;
        RECT 226.580 86.135 226.870 87.300 ;
        RECT 227.040 86.865 232.385 87.300 ;
        RECT 232.560 86.865 237.905 87.300 ;
        RECT 238.080 86.865 243.425 87.300 ;
        RECT 244.100 86.960 245.240 87.130 ;
        RECT 214.160 84.750 219.505 85.295 ;
        RECT 219.680 84.750 225.025 85.295 ;
        RECT 225.200 84.750 226.410 85.500 ;
        RECT 226.580 84.750 226.870 85.475 ;
        RECT 228.625 85.295 228.965 86.125 ;
        RECT 230.445 85.615 230.795 86.865 ;
        RECT 234.145 85.295 234.485 86.125 ;
        RECT 235.965 85.615 236.315 86.865 ;
        RECT 239.665 85.295 240.005 86.125 ;
        RECT 241.485 85.615 241.835 86.865 ;
        RECT 244.100 86.500 244.400 86.960 ;
        RECT 244.570 86.330 244.900 86.790 ;
        RECT 244.140 86.110 244.900 86.330 ;
        RECT 245.070 86.330 245.240 86.960 ;
        RECT 245.410 86.500 245.740 87.300 ;
        RECT 245.910 86.330 246.185 87.130 ;
        RECT 247.365 86.680 247.540 87.130 ;
        RECT 247.710 86.860 248.040 87.300 ;
        RECT 248.345 86.710 248.515 87.130 ;
        RECT 248.750 86.890 249.420 87.300 ;
        RECT 249.635 86.710 249.805 87.130 ;
        RECT 250.005 86.890 250.335 87.300 ;
        RECT 247.365 86.510 247.995 86.680 ;
        RECT 245.070 86.120 246.185 86.330 ;
        RECT 244.140 85.570 244.355 86.110 ;
        RECT 244.525 85.740 245.295 85.940 ;
        RECT 245.465 85.740 246.185 85.940 ;
        RECT 247.280 85.660 247.645 86.340 ;
        RECT 247.825 85.990 247.995 86.510 ;
        RECT 248.345 86.540 250.360 86.710 ;
        RECT 247.825 85.660 248.175 85.990 ;
        RECT 244.140 85.400 245.740 85.570 ;
        RECT 244.570 85.390 245.740 85.400 ;
        RECT 227.040 84.750 232.385 85.295 ;
        RECT 232.560 84.750 237.905 85.295 ;
        RECT 238.080 84.750 243.425 85.295 ;
        RECT 244.110 84.750 244.400 85.220 ;
        RECT 244.570 84.920 244.900 85.390 ;
        RECT 245.070 84.750 245.240 85.220 ;
        RECT 245.410 84.920 245.740 85.390 ;
        RECT 245.910 84.750 246.185 85.570 ;
        RECT 247.825 85.490 247.995 85.660 ;
        RECT 247.365 85.320 247.995 85.490 ;
        RECT 247.365 84.920 247.540 85.320 ;
        RECT 248.345 85.250 248.515 86.540 ;
        RECT 247.710 84.750 248.040 85.130 ;
        RECT 248.285 84.920 248.515 85.250 ;
        RECT 248.715 85.085 248.995 86.360 ;
        RECT 249.220 85.940 249.490 86.360 ;
        RECT 249.180 85.770 249.490 85.940 ;
        RECT 249.220 85.085 249.490 85.770 ;
        RECT 249.680 85.330 250.020 86.360 ;
        RECT 250.190 85.990 250.360 86.540 ;
        RECT 250.530 86.160 250.790 87.130 ;
        RECT 250.960 86.210 252.170 87.300 ;
        RECT 250.190 85.660 250.450 85.990 ;
        RECT 250.620 85.470 250.790 86.160 ;
        RECT 249.950 84.750 250.280 85.130 ;
        RECT 250.450 85.005 250.790 85.470 ;
        RECT 250.960 85.500 251.480 86.040 ;
        RECT 251.650 85.670 252.170 86.210 ;
        RECT 252.340 86.135 252.630 87.300 ;
        RECT 252.800 86.865 258.145 87.300 ;
        RECT 258.320 86.865 263.665 87.300 ;
        RECT 250.450 84.960 250.785 85.005 ;
        RECT 250.960 84.750 252.170 85.500 ;
        RECT 252.340 84.750 252.630 85.475 ;
        RECT 254.385 85.295 254.725 86.125 ;
        RECT 256.205 85.615 256.555 86.865 ;
        RECT 259.905 85.295 260.245 86.125 ;
        RECT 261.725 85.615 262.075 86.865 ;
        RECT 263.840 86.210 267.350 87.300 ;
        RECT 268.690 86.570 268.985 87.300 ;
        RECT 269.155 86.400 269.415 87.125 ;
        RECT 269.585 86.570 269.845 87.300 ;
        RECT 270.015 86.400 270.275 87.125 ;
        RECT 270.445 86.570 270.705 87.300 ;
        RECT 270.875 86.400 271.135 87.125 ;
        RECT 271.305 86.570 271.565 87.300 ;
        RECT 271.735 86.400 271.995 87.125 ;
        RECT 263.840 85.520 265.490 86.040 ;
        RECT 265.660 85.690 267.350 86.210 ;
        RECT 268.685 86.160 271.995 86.400 ;
        RECT 272.165 86.190 272.425 87.300 ;
        RECT 268.685 85.570 269.655 86.160 ;
        RECT 272.595 85.990 272.845 87.125 ;
        RECT 273.025 86.190 273.320 87.300 ;
        RECT 273.500 86.210 277.010 87.300 ;
        RECT 269.825 85.740 272.845 85.990 ;
        RECT 252.800 84.750 258.145 85.295 ;
        RECT 258.320 84.750 263.665 85.295 ;
        RECT 263.840 84.750 267.350 85.520 ;
        RECT 268.685 85.400 271.995 85.570 ;
        RECT 268.685 84.750 268.985 85.230 ;
        RECT 269.155 84.945 269.415 85.400 ;
        RECT 269.585 84.750 269.845 85.230 ;
        RECT 270.015 84.945 270.275 85.400 ;
        RECT 270.445 84.750 270.705 85.230 ;
        RECT 270.875 84.945 271.135 85.400 ;
        RECT 271.305 84.750 271.565 85.230 ;
        RECT 271.735 84.945 271.995 85.400 ;
        RECT 272.165 84.750 272.425 85.275 ;
        RECT 272.595 84.930 272.845 85.740 ;
        RECT 273.015 85.380 273.330 85.990 ;
        RECT 273.500 85.520 275.150 86.040 ;
        RECT 275.320 85.690 277.010 86.210 ;
        RECT 278.100 86.135 278.390 87.300 ;
        RECT 278.560 86.210 281.150 87.300 ;
        RECT 282.030 86.570 282.325 87.300 ;
        RECT 282.495 86.400 282.755 87.125 ;
        RECT 282.925 86.570 283.185 87.300 ;
        RECT 283.355 86.400 283.615 87.125 ;
        RECT 283.785 86.570 284.045 87.300 ;
        RECT 284.215 86.400 284.475 87.125 ;
        RECT 284.645 86.570 284.905 87.300 ;
        RECT 285.075 86.400 285.335 87.125 ;
        RECT 278.560 85.520 279.770 86.040 ;
        RECT 279.940 85.690 281.150 86.210 ;
        RECT 282.025 86.160 285.335 86.400 ;
        RECT 285.505 86.190 285.765 87.300 ;
        RECT 282.025 85.570 282.995 86.160 ;
        RECT 285.935 85.990 286.185 87.125 ;
        RECT 286.365 86.190 286.660 87.300 ;
        RECT 283.165 85.740 286.185 85.990 ;
        RECT 273.025 84.750 273.270 85.210 ;
        RECT 273.500 84.750 277.010 85.520 ;
        RECT 278.100 84.750 278.390 85.475 ;
        RECT 278.560 84.750 281.150 85.520 ;
        RECT 282.025 85.400 285.335 85.570 ;
        RECT 282.025 84.750 282.325 85.230 ;
        RECT 282.495 84.945 282.755 85.400 ;
        RECT 282.925 84.750 283.185 85.230 ;
        RECT 283.355 84.945 283.615 85.400 ;
        RECT 283.785 84.750 284.045 85.230 ;
        RECT 284.215 84.945 284.475 85.400 ;
        RECT 284.645 84.750 284.905 85.230 ;
        RECT 285.075 84.945 285.335 85.400 ;
        RECT 285.505 84.750 285.765 85.275 ;
        RECT 285.935 84.930 286.185 85.740 ;
        RECT 286.355 85.380 286.670 85.990 ;
        RECT 286.365 84.750 286.610 85.210 ;
        RECT 286.850 84.930 287.110 87.120 ;
        RECT 287.280 86.570 287.620 87.300 ;
        RECT 287.800 86.390 288.070 87.120 ;
        RECT 287.300 86.170 288.070 86.390 ;
        RECT 288.250 86.410 288.480 87.120 ;
        RECT 288.650 86.590 288.980 87.300 ;
        RECT 289.150 86.410 289.410 87.120 ;
        RECT 288.250 86.170 289.410 86.410 ;
        RECT 289.600 86.210 293.110 87.300 ;
        RECT 293.280 86.210 294.490 87.300 ;
        RECT 294.665 86.630 294.920 87.130 ;
        RECT 295.090 86.800 295.420 87.300 ;
        RECT 294.665 86.460 295.415 86.630 ;
        RECT 287.300 85.500 287.590 86.170 ;
        RECT 287.770 85.680 288.235 85.990 ;
        RECT 288.415 85.680 288.940 85.990 ;
        RECT 287.300 85.300 288.530 85.500 ;
        RECT 287.370 84.750 288.040 85.120 ;
        RECT 288.220 84.930 288.530 85.300 ;
        RECT 288.710 85.040 288.940 85.680 ;
        RECT 289.120 85.660 289.420 85.990 ;
        RECT 289.600 85.520 291.250 86.040 ;
        RECT 291.420 85.690 293.110 86.210 ;
        RECT 289.120 84.750 289.410 85.480 ;
        RECT 289.600 84.750 293.110 85.520 ;
        RECT 293.280 85.500 293.800 86.040 ;
        RECT 293.970 85.670 294.490 86.210 ;
        RECT 294.665 85.640 295.015 86.290 ;
        RECT 293.280 84.750 294.490 85.500 ;
        RECT 295.185 85.470 295.415 86.460 ;
        RECT 294.665 85.300 295.415 85.470 ;
        RECT 294.665 85.010 294.920 85.300 ;
        RECT 295.090 84.750 295.420 85.130 ;
        RECT 295.590 85.010 295.760 87.130 ;
        RECT 295.930 86.330 296.255 87.115 ;
        RECT 296.425 86.840 296.675 87.300 ;
        RECT 296.845 86.800 297.095 87.130 ;
        RECT 297.310 86.800 297.990 87.130 ;
        RECT 296.845 86.670 297.015 86.800 ;
        RECT 296.620 86.500 297.015 86.670 ;
        RECT 295.990 85.280 296.450 86.330 ;
        RECT 296.620 85.140 296.790 86.500 ;
        RECT 297.185 86.240 297.650 86.630 ;
        RECT 296.960 85.430 297.310 86.050 ;
        RECT 297.480 85.650 297.650 86.240 ;
        RECT 297.820 86.020 297.990 86.800 ;
        RECT 298.160 86.700 298.330 87.040 ;
        RECT 298.565 86.870 298.895 87.300 ;
        RECT 299.065 86.700 299.235 87.040 ;
        RECT 299.530 86.840 299.900 87.300 ;
        RECT 298.160 86.530 299.235 86.700 ;
        RECT 300.070 86.670 300.240 87.130 ;
        RECT 300.475 86.790 301.345 87.130 ;
        RECT 301.515 86.840 301.765 87.300 ;
        RECT 299.680 86.500 300.240 86.670 ;
        RECT 299.680 86.360 299.850 86.500 ;
        RECT 298.350 86.190 299.850 86.360 ;
        RECT 300.545 86.330 301.005 86.620 ;
        RECT 297.820 85.850 299.510 86.020 ;
        RECT 297.480 85.430 297.835 85.650 ;
        RECT 298.005 85.140 298.175 85.850 ;
        RECT 298.380 85.430 299.170 85.680 ;
        RECT 299.340 85.670 299.510 85.850 ;
        RECT 299.680 85.500 299.850 86.190 ;
        RECT 296.120 84.750 296.450 85.110 ;
        RECT 296.620 84.970 297.115 85.140 ;
        RECT 297.320 84.970 298.175 85.140 ;
        RECT 299.050 84.750 299.380 85.210 ;
        RECT 299.590 85.110 299.850 85.500 ;
        RECT 300.040 86.320 301.005 86.330 ;
        RECT 301.175 86.410 301.345 86.790 ;
        RECT 301.935 86.750 302.105 87.040 ;
        RECT 302.285 86.920 302.615 87.300 ;
        RECT 301.935 86.580 302.735 86.750 ;
        RECT 300.040 86.160 300.715 86.320 ;
        RECT 301.175 86.240 302.395 86.410 ;
        RECT 300.040 85.370 300.250 86.160 ;
        RECT 301.175 86.150 301.345 86.240 ;
        RECT 300.420 85.370 300.770 85.990 ;
        RECT 300.940 85.980 301.345 86.150 ;
        RECT 300.940 85.200 301.110 85.980 ;
        RECT 301.280 85.530 301.500 85.810 ;
        RECT 301.680 85.700 302.220 86.070 ;
        RECT 302.565 85.990 302.735 86.580 ;
        RECT 302.955 86.160 303.260 87.300 ;
        RECT 303.430 86.110 303.685 86.990 ;
        RECT 303.860 86.135 304.150 87.300 ;
        RECT 304.320 86.210 305.990 87.300 ;
        RECT 302.565 85.960 303.305 85.990 ;
        RECT 301.280 85.360 301.810 85.530 ;
        RECT 299.590 84.940 299.940 85.110 ;
        RECT 300.160 84.920 301.110 85.200 ;
        RECT 301.280 84.750 301.470 85.190 ;
        RECT 301.640 85.130 301.810 85.360 ;
        RECT 301.980 85.300 302.220 85.700 ;
        RECT 302.390 85.660 303.305 85.960 ;
        RECT 302.390 85.485 302.715 85.660 ;
        RECT 302.390 85.130 302.710 85.485 ;
        RECT 303.475 85.460 303.685 86.110 ;
        RECT 304.320 85.520 305.070 86.040 ;
        RECT 305.240 85.690 305.990 86.210 ;
        RECT 306.620 86.225 306.890 87.130 ;
        RECT 307.060 86.540 307.390 87.300 ;
        RECT 307.570 86.370 307.740 87.130 ;
        RECT 301.640 84.960 302.710 85.130 ;
        RECT 302.955 84.750 303.260 85.210 ;
        RECT 303.430 84.930 303.685 85.460 ;
        RECT 303.860 84.750 304.150 85.475 ;
        RECT 304.320 84.750 305.990 85.520 ;
        RECT 306.620 85.425 306.790 86.225 ;
        RECT 307.075 86.200 307.740 86.370 ;
        RECT 308.090 86.370 308.260 87.130 ;
        RECT 308.475 86.540 308.805 87.300 ;
        RECT 308.090 86.200 308.805 86.370 ;
        RECT 308.975 86.225 309.230 87.130 ;
        RECT 307.075 86.055 307.245 86.200 ;
        RECT 306.960 85.725 307.245 86.055 ;
        RECT 307.075 85.470 307.245 85.725 ;
        RECT 307.480 85.650 307.810 86.020 ;
        RECT 308.000 85.650 308.355 86.020 ;
        RECT 308.635 85.990 308.805 86.200 ;
        RECT 308.635 85.660 308.890 85.990 ;
        RECT 308.635 85.470 308.805 85.660 ;
        RECT 309.060 85.495 309.230 86.225 ;
        RECT 309.405 86.150 309.665 87.300 ;
        RECT 309.840 86.210 311.050 87.300 ;
        RECT 309.840 85.670 310.360 86.210 ;
        RECT 306.620 84.920 306.880 85.425 ;
        RECT 307.075 85.300 307.740 85.470 ;
        RECT 307.060 84.750 307.390 85.130 ;
        RECT 307.570 84.920 307.740 85.300 ;
        RECT 308.090 85.300 308.805 85.470 ;
        RECT 308.090 84.920 308.260 85.300 ;
        RECT 308.475 84.750 308.805 85.130 ;
        RECT 308.975 84.920 309.230 85.495 ;
        RECT 309.405 84.750 309.665 85.590 ;
        RECT 310.530 85.500 311.050 86.040 ;
        RECT 309.840 84.750 311.050 85.500 ;
        RECT 162.095 84.580 311.135 84.750 ;
        RECT 162.180 83.830 163.390 84.580 ;
        RECT 162.180 83.290 162.700 83.830 ;
        RECT 163.560 83.810 166.150 84.580 ;
        RECT 166.785 84.030 167.040 84.320 ;
        RECT 167.210 84.200 167.540 84.580 ;
        RECT 166.785 83.860 167.535 84.030 ;
        RECT 162.870 83.120 163.390 83.660 ;
        RECT 163.560 83.290 164.770 83.810 ;
        RECT 164.940 83.120 166.150 83.640 ;
        RECT 162.180 82.030 163.390 83.120 ;
        RECT 163.560 82.030 166.150 83.120 ;
        RECT 166.785 83.040 167.135 83.690 ;
        RECT 167.305 82.870 167.535 83.860 ;
        RECT 166.785 82.700 167.535 82.870 ;
        RECT 166.785 82.200 167.040 82.700 ;
        RECT 167.210 82.030 167.540 82.530 ;
        RECT 167.710 82.200 167.880 84.320 ;
        RECT 168.240 84.220 168.570 84.580 ;
        RECT 168.740 84.190 169.235 84.360 ;
        RECT 169.440 84.190 170.295 84.360 ;
        RECT 168.110 83.000 168.570 84.050 ;
        RECT 168.050 82.215 168.375 83.000 ;
        RECT 168.740 82.830 168.910 84.190 ;
        RECT 169.080 83.280 169.430 83.900 ;
        RECT 169.600 83.680 169.955 83.900 ;
        RECT 169.600 83.090 169.770 83.680 ;
        RECT 170.125 83.480 170.295 84.190 ;
        RECT 171.170 84.120 171.500 84.580 ;
        RECT 171.710 84.220 172.060 84.390 ;
        RECT 170.500 83.650 171.290 83.900 ;
        RECT 171.710 83.830 171.970 84.220 ;
        RECT 172.280 84.130 173.230 84.410 ;
        RECT 173.400 84.140 173.590 84.580 ;
        RECT 173.760 84.200 174.830 84.370 ;
        RECT 171.460 83.480 171.630 83.660 ;
        RECT 168.740 82.660 169.135 82.830 ;
        RECT 169.305 82.700 169.770 83.090 ;
        RECT 169.940 83.310 171.630 83.480 ;
        RECT 168.965 82.530 169.135 82.660 ;
        RECT 169.940 82.530 170.110 83.310 ;
        RECT 171.800 83.140 171.970 83.830 ;
        RECT 170.470 82.970 171.970 83.140 ;
        RECT 172.160 83.170 172.370 83.960 ;
        RECT 172.540 83.340 172.890 83.960 ;
        RECT 173.060 83.350 173.230 84.130 ;
        RECT 173.760 83.970 173.930 84.200 ;
        RECT 173.400 83.800 173.930 83.970 ;
        RECT 173.400 83.520 173.620 83.800 ;
        RECT 174.100 83.630 174.340 84.030 ;
        RECT 173.060 83.180 173.465 83.350 ;
        RECT 173.800 83.260 174.340 83.630 ;
        RECT 174.510 83.845 174.830 84.200 ;
        RECT 175.075 84.120 175.380 84.580 ;
        RECT 175.550 83.870 175.805 84.400 ;
        RECT 175.980 84.035 181.325 84.580 ;
        RECT 174.510 83.670 174.835 83.845 ;
        RECT 174.510 83.370 175.425 83.670 ;
        RECT 174.685 83.340 175.425 83.370 ;
        RECT 172.160 83.010 172.835 83.170 ;
        RECT 173.295 83.090 173.465 83.180 ;
        RECT 172.160 83.000 173.125 83.010 ;
        RECT 171.800 82.830 171.970 82.970 ;
        RECT 168.545 82.030 168.795 82.490 ;
        RECT 168.965 82.200 169.215 82.530 ;
        RECT 169.430 82.200 170.110 82.530 ;
        RECT 170.280 82.630 171.355 82.800 ;
        RECT 171.800 82.660 172.360 82.830 ;
        RECT 172.665 82.710 173.125 83.000 ;
        RECT 173.295 82.920 174.515 83.090 ;
        RECT 170.280 82.290 170.450 82.630 ;
        RECT 170.685 82.030 171.015 82.460 ;
        RECT 171.185 82.290 171.355 82.630 ;
        RECT 171.650 82.030 172.020 82.490 ;
        RECT 172.190 82.200 172.360 82.660 ;
        RECT 173.295 82.540 173.465 82.920 ;
        RECT 174.685 82.750 174.855 83.340 ;
        RECT 175.595 83.220 175.805 83.870 ;
        RECT 172.595 82.200 173.465 82.540 ;
        RECT 174.055 82.580 174.855 82.750 ;
        RECT 173.635 82.030 173.885 82.490 ;
        RECT 174.055 82.290 174.225 82.580 ;
        RECT 174.405 82.030 174.735 82.410 ;
        RECT 175.075 82.030 175.380 83.170 ;
        RECT 175.550 82.340 175.805 83.220 ;
        RECT 177.565 83.205 177.905 84.035 ;
        RECT 181.500 83.810 184.090 84.580 ;
        RECT 179.385 82.465 179.735 83.715 ;
        RECT 181.500 83.290 182.710 83.810 ;
        RECT 184.260 83.780 184.550 84.580 ;
        RECT 184.720 84.120 185.270 84.410 ;
        RECT 185.440 84.120 185.690 84.580 ;
        RECT 182.880 83.120 184.090 83.640 ;
        RECT 175.980 82.030 181.325 82.465 ;
        RECT 181.500 82.030 184.090 83.120 ;
        RECT 184.260 82.030 184.550 83.170 ;
        RECT 184.720 82.750 184.970 84.120 ;
        RECT 186.320 83.950 186.650 84.310 ;
        RECT 185.260 83.760 186.650 83.950 ;
        RECT 187.940 83.855 188.230 84.580 ;
        RECT 188.400 83.780 188.690 84.580 ;
        RECT 188.860 84.120 189.410 84.410 ;
        RECT 189.580 84.120 189.830 84.580 ;
        RECT 185.260 83.670 185.430 83.760 ;
        RECT 185.140 83.340 185.430 83.670 ;
        RECT 185.600 83.340 185.930 83.590 ;
        RECT 186.160 83.340 186.850 83.590 ;
        RECT 185.260 83.090 185.430 83.340 ;
        RECT 185.260 82.920 186.200 83.090 ;
        RECT 184.720 82.200 185.170 82.750 ;
        RECT 185.360 82.030 185.690 82.750 ;
        RECT 185.900 82.370 186.200 82.920 ;
        RECT 186.535 82.900 186.850 83.340 ;
        RECT 186.370 82.030 186.650 82.700 ;
        RECT 187.940 82.030 188.230 83.195 ;
        RECT 188.400 82.030 188.690 83.170 ;
        RECT 188.860 82.750 189.110 84.120 ;
        RECT 190.460 83.950 190.790 84.310 ;
        RECT 189.400 83.760 190.790 83.950 ;
        RECT 191.160 83.810 192.830 84.580 ;
        RECT 193.010 84.090 193.340 84.580 ;
        RECT 193.510 83.985 194.130 84.410 ;
        RECT 189.400 83.670 189.570 83.760 ;
        RECT 189.280 83.340 189.570 83.670 ;
        RECT 189.740 83.340 190.070 83.590 ;
        RECT 190.300 83.340 190.990 83.590 ;
        RECT 189.400 83.090 189.570 83.340 ;
        RECT 189.400 82.920 190.340 83.090 ;
        RECT 188.860 82.200 189.310 82.750 ;
        RECT 189.500 82.030 189.830 82.750 ;
        RECT 190.040 82.370 190.340 82.920 ;
        RECT 190.675 82.900 190.990 83.340 ;
        RECT 191.160 83.290 191.910 83.810 ;
        RECT 192.080 83.120 192.830 83.640 ;
        RECT 193.000 83.340 193.340 83.920 ;
        RECT 193.510 83.650 193.870 83.985 ;
        RECT 194.590 83.890 194.920 84.580 ;
        RECT 196.005 84.100 196.305 84.580 ;
        RECT 196.475 83.930 196.735 84.385 ;
        RECT 196.905 84.100 197.165 84.580 ;
        RECT 197.335 83.930 197.595 84.385 ;
        RECT 197.765 84.100 198.025 84.580 ;
        RECT 198.195 83.930 198.455 84.385 ;
        RECT 198.625 84.100 198.885 84.580 ;
        RECT 199.055 83.930 199.315 84.385 ;
        RECT 199.485 84.055 199.745 84.580 ;
        RECT 196.005 83.760 199.315 83.930 ;
        RECT 193.510 83.370 194.930 83.650 ;
        RECT 190.510 82.030 190.790 82.700 ;
        RECT 191.160 82.030 192.830 83.120 ;
        RECT 193.010 82.030 193.340 83.170 ;
        RECT 193.510 82.200 193.870 83.370 ;
        RECT 194.070 82.030 194.400 83.200 ;
        RECT 194.600 82.200 194.930 83.370 ;
        RECT 195.130 82.030 195.460 83.200 ;
        RECT 196.005 83.170 196.975 83.760 ;
        RECT 199.915 83.590 200.165 84.400 ;
        RECT 200.345 84.120 200.590 84.580 ;
        RECT 197.145 83.340 200.165 83.590 ;
        RECT 200.335 83.340 200.650 83.950 ;
        RECT 200.820 83.810 204.330 84.580 ;
        RECT 204.500 83.830 205.710 84.580 ;
        RECT 205.890 84.090 206.220 84.580 ;
        RECT 206.390 83.985 207.010 84.410 ;
        RECT 196.005 82.930 199.315 83.170 ;
        RECT 196.010 82.030 196.305 82.760 ;
        RECT 196.475 82.205 196.735 82.930 ;
        RECT 196.905 82.030 197.165 82.760 ;
        RECT 197.335 82.205 197.595 82.930 ;
        RECT 197.765 82.030 198.025 82.760 ;
        RECT 198.195 82.205 198.455 82.930 ;
        RECT 198.625 82.030 198.885 82.760 ;
        RECT 199.055 82.205 199.315 82.930 ;
        RECT 199.485 82.030 199.745 83.140 ;
        RECT 199.915 82.205 200.165 83.340 ;
        RECT 200.820 83.290 202.470 83.810 ;
        RECT 200.345 82.030 200.640 83.140 ;
        RECT 202.640 83.120 204.330 83.640 ;
        RECT 204.500 83.290 205.020 83.830 ;
        RECT 205.190 83.120 205.710 83.660 ;
        RECT 205.880 83.340 206.220 83.920 ;
        RECT 206.390 83.650 206.750 83.985 ;
        RECT 207.470 83.890 207.800 84.580 ;
        RECT 208.700 84.120 208.945 84.580 ;
        RECT 206.390 83.370 207.810 83.650 ;
        RECT 200.820 82.030 204.330 83.120 ;
        RECT 204.500 82.030 205.710 83.120 ;
        RECT 205.890 82.030 206.220 83.170 ;
        RECT 206.390 82.200 206.750 83.370 ;
        RECT 206.950 82.030 207.280 83.200 ;
        RECT 207.480 82.200 207.810 83.370 ;
        RECT 208.640 83.340 208.955 83.950 ;
        RECT 209.125 83.590 209.375 84.400 ;
        RECT 209.545 84.055 209.805 84.580 ;
        RECT 209.975 83.930 210.235 84.385 ;
        RECT 210.405 84.100 210.665 84.580 ;
        RECT 210.835 83.930 211.095 84.385 ;
        RECT 211.265 84.100 211.525 84.580 ;
        RECT 211.695 83.930 211.955 84.385 ;
        RECT 212.125 84.100 212.385 84.580 ;
        RECT 212.555 83.930 212.815 84.385 ;
        RECT 212.985 84.100 213.285 84.580 ;
        RECT 209.975 83.760 213.285 83.930 ;
        RECT 213.700 83.855 213.990 84.580 ;
        RECT 214.365 83.800 214.865 84.410 ;
        RECT 209.125 83.340 212.145 83.590 ;
        RECT 208.010 82.030 208.340 83.200 ;
        RECT 208.650 82.030 208.945 83.140 ;
        RECT 209.125 82.205 209.375 83.340 ;
        RECT 212.315 83.170 213.285 83.760 ;
        RECT 214.160 83.340 214.510 83.590 ;
        RECT 209.545 82.030 209.805 83.140 ;
        RECT 209.975 82.930 213.285 83.170 ;
        RECT 209.975 82.205 210.235 82.930 ;
        RECT 210.405 82.030 210.665 82.760 ;
        RECT 210.835 82.205 211.095 82.930 ;
        RECT 211.265 82.030 211.525 82.760 ;
        RECT 211.695 82.205 211.955 82.930 ;
        RECT 212.125 82.030 212.385 82.760 ;
        RECT 212.555 82.205 212.815 82.930 ;
        RECT 212.985 82.030 213.280 82.760 ;
        RECT 213.700 82.030 213.990 83.195 ;
        RECT 214.695 83.170 214.865 83.800 ;
        RECT 215.495 83.930 215.825 84.410 ;
        RECT 215.995 84.120 216.220 84.580 ;
        RECT 216.390 83.930 216.720 84.410 ;
        RECT 215.495 83.760 216.720 83.930 ;
        RECT 216.910 83.780 217.160 84.580 ;
        RECT 217.330 83.780 217.670 84.410 ;
        RECT 217.840 84.035 223.185 84.580 ;
        RECT 215.035 83.390 215.365 83.590 ;
        RECT 215.535 83.390 215.865 83.590 ;
        RECT 216.035 83.390 216.455 83.590 ;
        RECT 216.630 83.420 217.325 83.590 ;
        RECT 216.630 83.170 216.800 83.420 ;
        RECT 217.495 83.220 217.670 83.780 ;
        RECT 217.440 83.170 217.670 83.220 ;
        RECT 219.425 83.205 219.765 84.035 ;
        RECT 223.360 83.810 226.870 84.580 ;
        RECT 227.045 83.815 227.500 84.580 ;
        RECT 227.775 84.200 229.075 84.410 ;
        RECT 229.330 84.220 229.660 84.580 ;
        RECT 228.905 84.050 229.075 84.200 ;
        RECT 229.830 84.080 230.090 84.410 ;
        RECT 214.365 83.000 216.800 83.170 ;
        RECT 214.365 82.200 214.695 83.000 ;
        RECT 214.865 82.030 215.195 82.830 ;
        RECT 215.495 82.200 215.825 83.000 ;
        RECT 216.470 82.030 216.720 82.830 ;
        RECT 216.990 82.030 217.160 83.170 ;
        RECT 217.330 82.200 217.670 83.170 ;
        RECT 221.245 82.465 221.595 83.715 ;
        RECT 223.360 83.290 225.010 83.810 ;
        RECT 225.180 83.120 226.870 83.640 ;
        RECT 227.975 83.590 228.195 83.990 ;
        RECT 227.040 83.390 227.530 83.590 ;
        RECT 227.720 83.380 228.195 83.590 ;
        RECT 228.440 83.590 228.650 83.990 ;
        RECT 228.905 83.925 229.660 84.050 ;
        RECT 228.905 83.880 229.750 83.925 ;
        RECT 229.480 83.760 229.750 83.880 ;
        RECT 228.440 83.380 228.770 83.590 ;
        RECT 228.940 83.320 229.350 83.625 ;
        RECT 217.840 82.030 223.185 82.465 ;
        RECT 223.360 82.030 226.870 83.120 ;
        RECT 227.045 83.150 228.220 83.210 ;
        RECT 229.580 83.185 229.750 83.760 ;
        RECT 229.550 83.150 229.750 83.185 ;
        RECT 227.045 83.040 229.750 83.150 ;
        RECT 227.045 82.420 227.300 83.040 ;
        RECT 227.890 82.980 229.690 83.040 ;
        RECT 227.890 82.950 228.220 82.980 ;
        RECT 229.920 82.880 230.090 84.080 ;
        RECT 230.260 84.035 235.605 84.580 ;
        RECT 231.845 83.205 232.185 84.035 ;
        RECT 235.780 83.810 239.290 84.580 ;
        RECT 239.460 83.855 239.750 84.580 ;
        RECT 240.910 84.180 241.240 84.580 ;
        RECT 241.410 84.010 241.580 84.280 ;
        RECT 241.750 84.180 242.080 84.580 ;
        RECT 242.250 84.010 242.505 84.280 ;
        RECT 227.550 82.780 227.735 82.870 ;
        RECT 228.325 82.780 229.160 82.790 ;
        RECT 227.550 82.580 229.160 82.780 ;
        RECT 227.550 82.540 227.780 82.580 ;
        RECT 227.045 82.200 227.380 82.420 ;
        RECT 228.385 82.030 228.740 82.410 ;
        RECT 228.910 82.200 229.160 82.580 ;
        RECT 229.410 82.030 229.660 82.810 ;
        RECT 229.830 82.200 230.090 82.880 ;
        RECT 233.665 82.465 234.015 83.715 ;
        RECT 235.780 83.290 237.430 83.810 ;
        RECT 237.600 83.120 239.290 83.640 ;
        RECT 230.260 82.030 235.605 82.465 ;
        RECT 235.780 82.030 239.290 83.120 ;
        RECT 239.460 82.030 239.750 83.195 ;
        RECT 240.840 83.000 241.110 84.010 ;
        RECT 241.280 83.840 242.505 84.010 ;
        RECT 242.700 84.080 242.955 84.410 ;
        RECT 243.170 84.100 243.500 84.580 ;
        RECT 243.670 84.160 245.205 84.410 ;
        RECT 242.700 84.000 242.885 84.080 ;
        RECT 241.280 83.170 241.450 83.840 ;
        RECT 241.620 83.340 242.000 83.670 ;
        RECT 242.170 83.340 242.505 83.670 ;
        RECT 241.280 83.000 241.595 83.170 ;
        RECT 240.845 82.030 241.160 82.830 ;
        RECT 241.425 82.540 241.595 83.000 ;
        RECT 241.765 82.660 242.000 83.340 ;
        RECT 241.360 82.385 241.595 82.540 ;
        RECT 242.170 82.385 242.505 83.170 ;
        RECT 241.360 82.370 242.505 82.385 ;
        RECT 241.425 82.215 242.505 82.370 ;
        RECT 242.700 82.870 242.870 84.000 ;
        RECT 243.670 83.930 243.840 84.160 ;
        RECT 243.040 83.760 243.840 83.930 ;
        RECT 243.040 83.210 243.210 83.760 ;
        RECT 244.020 83.590 244.305 83.990 ;
        RECT 243.440 83.390 243.805 83.590 ;
        RECT 243.975 83.390 244.305 83.590 ;
        RECT 244.575 83.590 244.855 83.990 ;
        RECT 245.035 83.930 245.205 84.160 ;
        RECT 245.430 84.100 245.760 84.580 ;
        RECT 245.930 83.930 246.100 84.410 ;
        RECT 245.035 83.760 246.100 83.930 ;
        RECT 246.360 84.120 246.920 84.410 ;
        RECT 247.090 84.120 247.340 84.580 ;
        RECT 244.575 83.390 245.050 83.590 ;
        RECT 245.220 83.390 245.665 83.590 ;
        RECT 245.835 83.380 246.185 83.590 ;
        RECT 243.040 83.040 246.100 83.210 ;
        RECT 242.700 82.200 242.955 82.870 ;
        RECT 243.125 82.030 243.455 82.790 ;
        RECT 243.625 82.630 245.260 82.870 ;
        RECT 243.625 82.200 243.875 82.630 ;
        RECT 245.030 82.540 245.260 82.630 ;
        RECT 244.045 82.030 244.400 82.450 ;
        RECT 244.590 82.370 244.920 82.410 ;
        RECT 245.430 82.370 245.760 82.870 ;
        RECT 244.590 82.200 245.760 82.370 ;
        RECT 245.930 82.200 246.100 83.040 ;
        RECT 246.360 82.750 246.610 84.120 ;
        RECT 247.960 83.950 248.290 84.310 ;
        RECT 246.900 83.760 248.290 83.950 ;
        RECT 248.750 84.030 248.920 84.410 ;
        RECT 249.135 84.200 249.465 84.580 ;
        RECT 248.750 83.860 249.465 84.030 ;
        RECT 246.900 83.670 247.070 83.760 ;
        RECT 246.780 83.340 247.070 83.670 ;
        RECT 247.240 83.340 247.580 83.590 ;
        RECT 247.800 83.340 248.475 83.590 ;
        RECT 246.900 83.090 247.070 83.340 ;
        RECT 246.900 82.920 247.840 83.090 ;
        RECT 248.210 82.980 248.475 83.340 ;
        RECT 248.660 83.310 249.015 83.680 ;
        RECT 249.295 83.670 249.465 83.860 ;
        RECT 249.635 83.835 249.890 84.410 ;
        RECT 249.295 83.340 249.550 83.670 ;
        RECT 249.295 83.130 249.465 83.340 ;
        RECT 246.360 82.200 246.820 82.750 ;
        RECT 247.010 82.030 247.340 82.750 ;
        RECT 247.540 82.370 247.840 82.920 ;
        RECT 248.750 82.960 249.465 83.130 ;
        RECT 249.720 83.105 249.890 83.835 ;
        RECT 250.065 83.740 250.325 84.580 ;
        RECT 250.590 84.030 250.760 84.410 ;
        RECT 250.975 84.200 251.305 84.580 ;
        RECT 250.590 83.860 251.305 84.030 ;
        RECT 250.500 83.310 250.855 83.680 ;
        RECT 251.135 83.670 251.305 83.860 ;
        RECT 251.475 83.835 251.730 84.410 ;
        RECT 251.135 83.340 251.390 83.670 ;
        RECT 248.010 82.030 248.290 82.700 ;
        RECT 248.750 82.200 248.920 82.960 ;
        RECT 249.135 82.030 249.465 82.790 ;
        RECT 249.635 82.200 249.890 83.105 ;
        RECT 250.065 82.030 250.325 83.180 ;
        RECT 251.135 83.130 251.305 83.340 ;
        RECT 250.590 82.960 251.305 83.130 ;
        RECT 251.560 83.105 251.730 83.835 ;
        RECT 251.905 83.740 252.165 84.580 ;
        RECT 252.345 84.180 252.680 84.580 ;
        RECT 252.850 84.010 253.055 84.410 ;
        RECT 253.265 84.100 253.540 84.580 ;
        RECT 253.750 84.080 254.010 84.410 ;
        RECT 252.370 83.840 253.055 84.010 ;
        RECT 250.590 82.200 250.760 82.960 ;
        RECT 250.975 82.030 251.305 82.790 ;
        RECT 251.475 82.200 251.730 83.105 ;
        RECT 251.905 82.030 252.165 83.180 ;
        RECT 252.370 82.810 252.710 83.840 ;
        RECT 252.880 83.170 253.130 83.670 ;
        RECT 253.310 83.340 253.670 83.920 ;
        RECT 253.840 83.170 254.010 84.080 ;
        RECT 254.180 84.035 259.525 84.580 ;
        RECT 260.630 84.080 260.960 84.580 ;
        RECT 255.765 83.205 256.105 84.035 ;
        RECT 261.160 84.010 261.330 84.360 ;
        RECT 261.530 84.180 261.860 84.580 ;
        RECT 262.030 84.010 262.200 84.360 ;
        RECT 262.370 84.180 262.750 84.580 ;
        RECT 252.880 83.000 254.010 83.170 ;
        RECT 252.370 82.635 253.035 82.810 ;
        RECT 252.345 82.030 252.680 82.455 ;
        RECT 252.850 82.230 253.035 82.635 ;
        RECT 253.240 82.030 253.570 82.810 ;
        RECT 253.740 82.230 254.010 83.000 ;
        RECT 257.585 82.465 257.935 83.715 ;
        RECT 260.625 83.340 260.975 83.910 ;
        RECT 261.160 83.840 262.770 84.010 ;
        RECT 262.940 83.905 263.210 84.250 ;
        RECT 262.600 83.670 262.770 83.840 ;
        RECT 260.625 82.880 260.945 83.170 ;
        RECT 261.145 83.050 261.855 83.670 ;
        RECT 262.025 83.340 262.430 83.670 ;
        RECT 262.600 83.340 262.870 83.670 ;
        RECT 262.600 83.170 262.770 83.340 ;
        RECT 263.040 83.170 263.210 83.905 ;
        RECT 263.380 83.810 265.050 84.580 ;
        RECT 265.220 83.855 265.510 84.580 ;
        RECT 265.880 83.950 266.210 84.310 ;
        RECT 266.830 84.120 267.080 84.580 ;
        RECT 267.250 84.120 267.810 84.410 ;
        RECT 263.380 83.290 264.130 83.810 ;
        RECT 265.880 83.760 267.270 83.950 ;
        RECT 267.100 83.670 267.270 83.760 ;
        RECT 262.045 83.000 262.770 83.170 ;
        RECT 262.045 82.880 262.215 83.000 ;
        RECT 260.625 82.710 262.215 82.880 ;
        RECT 254.180 82.030 259.525 82.465 ;
        RECT 260.625 82.250 262.280 82.540 ;
        RECT 262.450 82.030 262.730 82.830 ;
        RECT 262.940 82.200 263.210 83.170 ;
        RECT 264.300 83.120 265.050 83.640 ;
        RECT 265.695 83.340 266.370 83.590 ;
        RECT 266.590 83.340 266.930 83.590 ;
        RECT 267.100 83.340 267.390 83.670 ;
        RECT 263.380 82.030 265.050 83.120 ;
        RECT 265.220 82.030 265.510 83.195 ;
        RECT 265.695 82.980 265.960 83.340 ;
        RECT 267.100 83.090 267.270 83.340 ;
        RECT 266.330 82.920 267.270 83.090 ;
        RECT 265.880 82.030 266.160 82.700 ;
        RECT 266.330 82.370 266.630 82.920 ;
        RECT 267.560 82.750 267.810 84.120 ;
        RECT 268.540 84.115 268.790 84.580 ;
        RECT 268.960 83.940 269.130 84.410 ;
        RECT 269.380 84.120 269.550 84.580 ;
        RECT 269.800 83.940 269.970 84.410 ;
        RECT 270.220 84.120 270.390 84.580 ;
        RECT 270.640 83.940 270.810 84.410 ;
        RECT 271.180 84.120 271.445 84.580 ;
        RECT 271.660 84.035 277.005 84.580 ;
        RECT 268.440 83.760 270.810 83.940 ;
        RECT 268.440 83.170 268.790 83.760 ;
        RECT 268.960 83.340 271.470 83.590 ;
        RECT 273.245 83.205 273.585 84.035 ;
        RECT 277.380 83.950 277.710 84.310 ;
        RECT 278.340 84.120 278.590 84.580 ;
        RECT 278.760 84.120 279.310 84.410 ;
        RECT 277.380 83.760 278.770 83.950 ;
        RECT 268.440 83.000 270.890 83.170 ;
        RECT 268.440 82.980 269.210 83.000 ;
        RECT 266.830 82.030 267.160 82.750 ;
        RECT 267.350 82.200 267.810 82.750 ;
        RECT 268.540 82.030 268.710 82.490 ;
        RECT 268.880 82.200 269.210 82.980 ;
        RECT 269.380 82.030 269.550 82.830 ;
        RECT 269.720 82.200 270.050 83.000 ;
        RECT 270.220 82.030 270.390 82.830 ;
        RECT 270.560 82.200 270.890 83.000 ;
        RECT 271.150 82.030 271.445 83.170 ;
        RECT 275.065 82.465 275.415 83.715 ;
        RECT 278.600 83.670 278.770 83.760 ;
        RECT 277.180 83.340 277.870 83.590 ;
        RECT 278.100 83.340 278.430 83.590 ;
        RECT 278.600 83.340 278.890 83.670 ;
        RECT 277.180 82.900 277.495 83.340 ;
        RECT 278.600 83.090 278.770 83.340 ;
        RECT 277.830 82.920 278.770 83.090 ;
        RECT 271.660 82.030 277.005 82.465 ;
        RECT 277.380 82.030 277.660 82.700 ;
        RECT 277.830 82.370 278.130 82.920 ;
        RECT 279.060 82.750 279.310 84.120 ;
        RECT 279.480 83.780 279.770 84.580 ;
        RECT 279.940 83.810 281.610 84.580 ;
        RECT 281.880 84.115 282.130 84.580 ;
        RECT 282.300 83.940 282.470 84.410 ;
        RECT 282.720 84.120 282.890 84.580 ;
        RECT 283.140 83.940 283.310 84.410 ;
        RECT 283.560 84.120 283.730 84.580 ;
        RECT 283.980 83.940 284.150 84.410 ;
        RECT 284.520 84.120 284.785 84.580 ;
        RECT 285.000 84.035 290.345 84.580 ;
        RECT 279.940 83.290 280.690 83.810 ;
        RECT 281.780 83.760 284.150 83.940 ;
        RECT 278.340 82.030 278.670 82.750 ;
        RECT 278.860 82.200 279.310 82.750 ;
        RECT 279.480 82.030 279.770 83.170 ;
        RECT 280.860 83.120 281.610 83.640 ;
        RECT 279.940 82.030 281.610 83.120 ;
        RECT 281.780 83.170 282.130 83.760 ;
        RECT 282.300 83.340 284.810 83.590 ;
        RECT 286.585 83.205 286.925 84.035 ;
        RECT 290.980 83.855 291.270 84.580 ;
        RECT 292.110 83.890 292.440 84.580 ;
        RECT 292.900 83.985 293.520 84.410 ;
        RECT 293.690 84.090 294.020 84.580 ;
        RECT 281.780 83.000 284.230 83.170 ;
        RECT 281.780 82.980 282.550 83.000 ;
        RECT 281.880 82.030 282.050 82.490 ;
        RECT 282.220 82.200 282.550 82.980 ;
        RECT 282.720 82.030 282.890 82.830 ;
        RECT 283.060 82.200 283.390 83.000 ;
        RECT 283.560 82.030 283.730 82.830 ;
        RECT 283.900 82.200 284.230 83.000 ;
        RECT 284.490 82.030 284.785 83.170 ;
        RECT 288.405 82.465 288.755 83.715 ;
        RECT 293.160 83.650 293.520 83.985 ;
        RECT 292.100 83.370 293.520 83.650 ;
        RECT 285.000 82.030 290.345 82.465 ;
        RECT 290.980 82.030 291.270 83.195 ;
        RECT 291.570 82.030 291.900 83.200 ;
        RECT 292.100 82.200 292.430 83.370 ;
        RECT 292.630 82.030 292.960 83.200 ;
        RECT 293.160 82.200 293.520 83.370 ;
        RECT 293.690 83.340 294.030 83.920 ;
        RECT 294.200 83.810 295.870 84.580 ;
        RECT 296.045 84.030 296.300 84.320 ;
        RECT 296.470 84.200 296.800 84.580 ;
        RECT 296.045 83.860 296.795 84.030 ;
        RECT 294.200 83.290 294.950 83.810 ;
        RECT 293.690 82.030 294.020 83.170 ;
        RECT 295.120 83.120 295.870 83.640 ;
        RECT 294.200 82.030 295.870 83.120 ;
        RECT 296.045 83.040 296.395 83.690 ;
        RECT 296.565 82.870 296.795 83.860 ;
        RECT 296.045 82.700 296.795 82.870 ;
        RECT 296.045 82.200 296.300 82.700 ;
        RECT 296.470 82.030 296.800 82.530 ;
        RECT 296.970 82.200 297.140 84.320 ;
        RECT 297.500 84.220 297.830 84.580 ;
        RECT 298.000 84.190 298.495 84.360 ;
        RECT 298.700 84.190 299.555 84.360 ;
        RECT 297.370 83.000 297.830 84.050 ;
        RECT 297.310 82.215 297.635 83.000 ;
        RECT 298.000 82.830 298.170 84.190 ;
        RECT 298.340 83.280 298.690 83.900 ;
        RECT 298.860 83.680 299.215 83.900 ;
        RECT 298.860 83.090 299.030 83.680 ;
        RECT 299.385 83.480 299.555 84.190 ;
        RECT 300.430 84.120 300.760 84.580 ;
        RECT 300.970 84.220 301.320 84.390 ;
        RECT 299.760 83.650 300.550 83.900 ;
        RECT 300.970 83.830 301.230 84.220 ;
        RECT 301.540 84.130 302.490 84.410 ;
        RECT 302.660 84.140 302.850 84.580 ;
        RECT 303.020 84.200 304.090 84.370 ;
        RECT 300.720 83.480 300.890 83.660 ;
        RECT 298.000 82.660 298.395 82.830 ;
        RECT 298.565 82.700 299.030 83.090 ;
        RECT 299.200 83.310 300.890 83.480 ;
        RECT 298.225 82.530 298.395 82.660 ;
        RECT 299.200 82.530 299.370 83.310 ;
        RECT 301.060 83.140 301.230 83.830 ;
        RECT 299.730 82.970 301.230 83.140 ;
        RECT 301.420 83.170 301.630 83.960 ;
        RECT 301.800 83.340 302.150 83.960 ;
        RECT 302.320 83.350 302.490 84.130 ;
        RECT 303.020 83.970 303.190 84.200 ;
        RECT 302.660 83.800 303.190 83.970 ;
        RECT 302.660 83.520 302.880 83.800 ;
        RECT 303.360 83.630 303.600 84.030 ;
        RECT 302.320 83.180 302.725 83.350 ;
        RECT 303.060 83.260 303.600 83.630 ;
        RECT 303.770 83.845 304.090 84.200 ;
        RECT 304.335 84.120 304.640 84.580 ;
        RECT 304.810 83.870 305.065 84.400 ;
        RECT 303.770 83.670 304.095 83.845 ;
        RECT 303.770 83.370 304.685 83.670 ;
        RECT 303.945 83.340 304.685 83.370 ;
        RECT 301.420 83.010 302.095 83.170 ;
        RECT 302.555 83.090 302.725 83.180 ;
        RECT 301.420 83.000 302.385 83.010 ;
        RECT 301.060 82.830 301.230 82.970 ;
        RECT 297.805 82.030 298.055 82.490 ;
        RECT 298.225 82.200 298.475 82.530 ;
        RECT 298.690 82.200 299.370 82.530 ;
        RECT 299.540 82.630 300.615 82.800 ;
        RECT 301.060 82.660 301.620 82.830 ;
        RECT 301.925 82.710 302.385 83.000 ;
        RECT 302.555 82.920 303.775 83.090 ;
        RECT 299.540 82.290 299.710 82.630 ;
        RECT 299.945 82.030 300.275 82.460 ;
        RECT 300.445 82.290 300.615 82.630 ;
        RECT 300.910 82.030 301.280 82.490 ;
        RECT 301.450 82.200 301.620 82.660 ;
        RECT 302.555 82.540 302.725 82.920 ;
        RECT 303.945 82.750 304.115 83.340 ;
        RECT 304.855 83.220 305.065 83.870 ;
        RECT 305.240 83.810 308.750 84.580 ;
        RECT 309.840 83.830 311.050 84.580 ;
        RECT 305.240 83.290 306.890 83.810 ;
        RECT 301.855 82.200 302.725 82.540 ;
        RECT 303.315 82.580 304.115 82.750 ;
        RECT 302.895 82.030 303.145 82.490 ;
        RECT 303.315 82.290 303.485 82.580 ;
        RECT 303.665 82.030 303.995 82.410 ;
        RECT 304.335 82.030 304.640 83.170 ;
        RECT 304.810 82.340 305.065 83.220 ;
        RECT 307.060 83.120 308.750 83.640 ;
        RECT 305.240 82.030 308.750 83.120 ;
        RECT 309.840 83.120 310.360 83.660 ;
        RECT 310.530 83.290 311.050 83.830 ;
        RECT 309.840 82.030 311.050 83.120 ;
        RECT 162.095 81.860 311.135 82.030 ;
        RECT 162.180 80.770 163.390 81.860 ;
        RECT 163.560 81.425 168.905 81.860 ;
        RECT 162.180 80.060 162.700 80.600 ;
        RECT 162.870 80.230 163.390 80.770 ;
        RECT 162.180 79.310 163.390 80.060 ;
        RECT 165.145 79.855 165.485 80.685 ;
        RECT 166.965 80.175 167.315 81.425 ;
        RECT 169.080 80.770 170.750 81.860 ;
        RECT 169.080 80.080 169.830 80.600 ;
        RECT 170.000 80.250 170.750 80.770 ;
        RECT 170.925 80.720 171.260 81.690 ;
        RECT 171.430 80.720 171.600 81.860 ;
        RECT 171.770 81.520 173.800 81.690 ;
        RECT 163.560 79.310 168.905 79.855 ;
        RECT 169.080 79.310 170.750 80.080 ;
        RECT 170.925 80.050 171.095 80.720 ;
        RECT 171.770 80.550 171.940 81.520 ;
        RECT 171.265 80.220 171.520 80.550 ;
        RECT 171.745 80.220 171.940 80.550 ;
        RECT 172.110 81.180 173.235 81.350 ;
        RECT 171.350 80.050 171.520 80.220 ;
        RECT 172.110 80.050 172.280 81.180 ;
        RECT 170.925 79.480 171.180 80.050 ;
        RECT 171.350 79.880 172.280 80.050 ;
        RECT 172.450 80.840 173.460 81.010 ;
        RECT 172.450 80.040 172.620 80.840 ;
        RECT 172.825 80.160 173.100 80.640 ;
        RECT 172.820 79.990 173.100 80.160 ;
        RECT 172.105 79.845 172.280 79.880 ;
        RECT 171.350 79.310 171.680 79.710 ;
        RECT 172.105 79.480 172.635 79.845 ;
        RECT 172.825 79.480 173.100 79.990 ;
        RECT 173.270 79.480 173.460 80.840 ;
        RECT 173.630 80.855 173.800 81.520 ;
        RECT 173.970 81.100 174.140 81.860 ;
        RECT 174.375 81.100 174.890 81.510 ;
        RECT 173.630 80.665 174.380 80.855 ;
        RECT 174.550 80.290 174.890 81.100 ;
        RECT 175.060 80.695 175.350 81.860 ;
        RECT 175.525 80.720 175.860 81.690 ;
        RECT 176.030 80.720 176.200 81.860 ;
        RECT 176.370 81.520 178.400 81.690 ;
        RECT 173.660 80.120 174.890 80.290 ;
        RECT 173.640 79.310 174.150 79.845 ;
        RECT 174.370 79.515 174.615 80.120 ;
        RECT 175.525 80.050 175.695 80.720 ;
        RECT 176.370 80.550 176.540 81.520 ;
        RECT 175.865 80.220 176.120 80.550 ;
        RECT 176.345 80.220 176.540 80.550 ;
        RECT 176.710 81.180 177.835 81.350 ;
        RECT 175.950 80.050 176.120 80.220 ;
        RECT 176.710 80.050 176.880 81.180 ;
        RECT 175.060 79.310 175.350 80.035 ;
        RECT 175.525 79.480 175.780 80.050 ;
        RECT 175.950 79.880 176.880 80.050 ;
        RECT 177.050 80.840 178.060 81.010 ;
        RECT 177.050 80.040 177.220 80.840 ;
        RECT 176.705 79.845 176.880 79.880 ;
        RECT 175.950 79.310 176.280 79.710 ;
        RECT 176.705 79.480 177.235 79.845 ;
        RECT 177.425 79.820 177.700 80.640 ;
        RECT 177.420 79.650 177.700 79.820 ;
        RECT 177.425 79.480 177.700 79.650 ;
        RECT 177.870 79.480 178.060 80.840 ;
        RECT 178.230 80.855 178.400 81.520 ;
        RECT 178.570 81.100 178.740 81.860 ;
        RECT 178.975 81.100 179.490 81.510 ;
        RECT 179.660 81.425 185.005 81.860 ;
        RECT 178.230 80.665 178.980 80.855 ;
        RECT 179.150 80.290 179.490 81.100 ;
        RECT 178.260 80.120 179.490 80.290 ;
        RECT 178.240 79.310 178.750 79.845 ;
        RECT 178.970 79.515 179.215 80.120 ;
        RECT 181.245 79.855 181.585 80.685 ;
        RECT 183.065 80.175 183.415 81.425 ;
        RECT 185.180 80.770 188.690 81.860 ;
        RECT 188.960 81.400 189.130 81.860 ;
        RECT 189.300 80.910 189.630 81.690 ;
        RECT 189.800 81.060 189.970 81.860 ;
        RECT 185.180 80.080 186.830 80.600 ;
        RECT 187.000 80.250 188.690 80.770 ;
        RECT 188.860 80.890 189.630 80.910 ;
        RECT 190.140 80.890 190.470 81.690 ;
        RECT 190.640 81.060 190.810 81.860 ;
        RECT 190.980 80.890 191.310 81.690 ;
        RECT 188.860 80.720 191.310 80.890 ;
        RECT 191.570 80.720 191.865 81.860 ;
        RECT 192.080 80.770 193.750 81.860 ;
        RECT 194.390 81.140 194.720 81.860 ;
        RECT 188.860 80.130 189.210 80.720 ;
        RECT 189.380 80.300 191.890 80.550 ;
        RECT 179.660 79.310 185.005 79.855 ;
        RECT 185.180 79.310 188.690 80.080 ;
        RECT 188.860 79.950 191.230 80.130 ;
        RECT 188.960 79.310 189.210 79.775 ;
        RECT 189.380 79.480 189.550 79.950 ;
        RECT 189.800 79.310 189.970 79.770 ;
        RECT 190.220 79.480 190.390 79.950 ;
        RECT 190.640 79.310 190.810 79.770 ;
        RECT 191.060 79.480 191.230 79.950 ;
        RECT 192.080 80.080 192.830 80.600 ;
        RECT 193.000 80.250 193.750 80.770 ;
        RECT 194.380 80.500 194.610 80.840 ;
        RECT 194.900 80.500 195.115 81.615 ;
        RECT 195.310 80.915 195.640 81.690 ;
        RECT 195.810 81.085 196.520 81.860 ;
        RECT 195.310 80.700 196.460 80.915 ;
        RECT 194.380 80.300 194.710 80.500 ;
        RECT 194.900 80.320 195.350 80.500 ;
        RECT 195.020 80.300 195.350 80.320 ;
        RECT 195.520 80.300 195.990 80.530 ;
        RECT 196.175 80.130 196.460 80.700 ;
        RECT 196.690 80.255 196.970 81.690 ;
        RECT 197.140 80.770 200.650 81.860 ;
        RECT 191.600 79.310 191.865 79.770 ;
        RECT 192.080 79.310 193.750 80.080 ;
        RECT 194.380 79.940 195.560 80.130 ;
        RECT 194.380 79.480 194.720 79.940 ;
        RECT 195.230 79.860 195.560 79.940 ;
        RECT 195.750 79.940 196.460 80.130 ;
        RECT 195.750 79.800 196.050 79.940 ;
        RECT 195.735 79.790 196.050 79.800 ;
        RECT 195.725 79.780 196.050 79.790 ;
        RECT 195.715 79.775 196.050 79.780 ;
        RECT 194.890 79.310 195.060 79.770 ;
        RECT 195.710 79.765 196.050 79.775 ;
        RECT 195.705 79.760 196.050 79.765 ;
        RECT 195.700 79.750 196.050 79.760 ;
        RECT 195.695 79.745 196.050 79.750 ;
        RECT 195.690 79.480 196.050 79.745 ;
        RECT 196.290 79.310 196.460 79.770 ;
        RECT 196.630 79.480 196.970 80.255 ;
        RECT 197.140 80.080 198.790 80.600 ;
        RECT 198.960 80.250 200.650 80.770 ;
        RECT 200.820 80.695 201.110 81.860 ;
        RECT 201.280 80.770 204.790 81.860 ;
        RECT 201.280 80.080 202.930 80.600 ;
        RECT 203.100 80.250 204.790 80.770 ;
        RECT 204.985 80.850 205.280 81.690 ;
        RECT 205.450 81.020 205.700 81.860 ;
        RECT 205.870 81.190 206.120 81.690 ;
        RECT 206.290 81.360 206.540 81.860 ;
        RECT 206.710 81.190 206.960 81.690 ;
        RECT 207.130 81.360 207.380 81.860 ;
        RECT 207.650 81.520 211.260 81.690 ;
        RECT 207.650 81.360 207.900 81.520 ;
        RECT 208.490 81.360 208.740 81.520 ;
        RECT 208.070 81.190 208.320 81.350 ;
        RECT 208.910 81.190 209.160 81.350 ;
        RECT 205.870 81.020 209.160 81.190 ;
        RECT 209.330 81.020 209.580 81.520 ;
        RECT 209.750 80.850 210.000 81.350 ;
        RECT 210.170 81.020 210.420 81.520 ;
        RECT 210.590 80.850 210.840 81.350 ;
        RECT 211.010 81.020 211.260 81.520 ;
        RECT 211.430 80.850 211.635 81.640 ;
        RECT 204.985 80.680 209.580 80.850 ;
        RECT 209.750 80.680 211.635 80.850 ;
        RECT 211.885 80.850 212.180 81.690 ;
        RECT 212.350 81.020 212.600 81.860 ;
        RECT 212.770 81.190 213.020 81.690 ;
        RECT 213.190 81.360 213.440 81.860 ;
        RECT 213.610 81.190 213.860 81.690 ;
        RECT 214.030 81.360 214.280 81.860 ;
        RECT 214.550 81.520 218.160 81.690 ;
        RECT 214.550 81.360 214.800 81.520 ;
        RECT 215.390 81.360 215.640 81.520 ;
        RECT 214.970 81.190 215.220 81.350 ;
        RECT 215.810 81.190 216.060 81.350 ;
        RECT 212.770 81.020 216.060 81.190 ;
        RECT 216.230 81.020 216.480 81.520 ;
        RECT 216.650 80.850 216.900 81.350 ;
        RECT 217.070 81.020 217.320 81.520 ;
        RECT 217.490 80.850 217.740 81.350 ;
        RECT 217.910 81.020 218.160 81.520 ;
        RECT 218.330 80.850 218.535 81.640 ;
        RECT 211.885 80.680 216.480 80.850 ;
        RECT 216.650 80.680 218.535 80.850 ;
        RECT 218.760 80.770 222.270 81.860 ;
        RECT 222.440 80.770 223.650 81.860 ;
        RECT 223.820 81.355 224.450 81.860 ;
        RECT 204.985 80.300 205.320 80.510 ;
        RECT 205.490 80.130 205.660 80.680 ;
        RECT 209.410 80.510 209.580 80.680 ;
        RECT 205.910 80.300 207.565 80.510 ;
        RECT 207.910 80.300 209.175 80.510 ;
        RECT 209.410 80.300 211.000 80.510 ;
        RECT 211.295 80.130 211.635 80.680 ;
        RECT 211.885 80.300 212.220 80.510 ;
        RECT 212.390 80.130 212.560 80.680 ;
        RECT 216.310 80.510 216.480 80.680 ;
        RECT 212.810 80.300 214.465 80.510 ;
        RECT 214.810 80.300 216.075 80.510 ;
        RECT 216.310 80.300 217.900 80.510 ;
        RECT 218.195 80.130 218.535 80.680 ;
        RECT 197.140 79.310 200.650 80.080 ;
        RECT 200.820 79.310 201.110 80.035 ;
        RECT 201.280 79.310 204.790 80.080 ;
        RECT 204.985 79.960 205.660 80.130 ;
        RECT 204.985 79.480 205.320 79.960 ;
        RECT 205.830 79.950 211.635 80.130 ;
        RECT 205.490 79.310 205.660 79.780 ;
        RECT 205.830 79.480 206.160 79.950 ;
        RECT 206.330 79.310 206.500 79.780 ;
        RECT 206.670 79.480 207.000 79.950 ;
        RECT 207.170 79.310 207.860 79.780 ;
        RECT 208.030 79.480 208.360 79.950 ;
        RECT 208.530 79.310 208.700 79.780 ;
        RECT 208.870 79.480 209.200 79.950 ;
        RECT 209.370 79.310 209.540 79.780 ;
        RECT 209.710 79.480 210.040 79.950 ;
        RECT 210.210 79.310 210.380 79.780 ;
        RECT 210.550 79.480 210.880 79.950 ;
        RECT 211.050 79.310 211.220 79.780 ;
        RECT 211.390 79.540 211.635 79.950 ;
        RECT 211.885 79.960 212.560 80.130 ;
        RECT 211.885 79.480 212.220 79.960 ;
        RECT 212.730 79.950 218.535 80.130 ;
        RECT 212.390 79.310 212.560 79.780 ;
        RECT 212.730 79.480 213.060 79.950 ;
        RECT 213.230 79.310 213.400 79.780 ;
        RECT 213.570 79.480 213.900 79.950 ;
        RECT 214.070 79.310 214.760 79.780 ;
        RECT 214.930 79.480 215.260 79.950 ;
        RECT 215.430 79.310 215.600 79.780 ;
        RECT 215.770 79.480 216.100 79.950 ;
        RECT 216.270 79.310 216.440 79.780 ;
        RECT 216.610 79.480 216.940 79.950 ;
        RECT 217.110 79.310 217.280 79.780 ;
        RECT 217.450 79.480 217.780 79.950 ;
        RECT 217.950 79.310 218.120 79.780 ;
        RECT 218.290 79.540 218.535 79.950 ;
        RECT 218.760 80.080 220.410 80.600 ;
        RECT 220.580 80.250 222.270 80.770 ;
        RECT 218.760 79.310 222.270 80.080 ;
        RECT 222.440 80.060 222.960 80.600 ;
        RECT 223.130 80.230 223.650 80.770 ;
        RECT 223.835 80.820 224.090 81.185 ;
        RECT 224.260 81.180 224.450 81.355 ;
        RECT 224.630 81.350 225.105 81.690 ;
        RECT 224.260 80.990 224.590 81.180 ;
        RECT 224.815 80.820 225.065 81.115 ;
        RECT 225.290 81.015 225.505 81.860 ;
        RECT 225.705 81.020 225.980 81.690 ;
        RECT 223.835 80.650 225.625 80.820 ;
        RECT 225.810 80.670 225.980 81.020 ;
        RECT 226.150 80.850 226.410 81.860 ;
        RECT 226.580 80.695 226.870 81.860 ;
        RECT 227.040 80.770 228.710 81.860 ;
        RECT 222.440 79.310 223.650 80.060 ;
        RECT 223.820 79.990 224.205 80.470 ;
        RECT 224.375 79.795 224.630 80.650 ;
        RECT 223.840 79.530 224.630 79.795 ;
        RECT 224.800 79.975 225.210 80.470 ;
        RECT 225.395 80.220 225.625 80.650 ;
        RECT 225.795 80.150 226.410 80.670 ;
        RECT 224.800 79.530 225.030 79.975 ;
        RECT 225.795 79.940 225.965 80.150 ;
        RECT 227.040 80.080 227.790 80.600 ;
        RECT 227.960 80.250 228.710 80.770 ;
        RECT 228.900 81.020 229.155 81.690 ;
        RECT 229.325 81.100 229.655 81.860 ;
        RECT 229.825 81.260 230.075 81.690 ;
        RECT 230.245 81.440 230.600 81.860 ;
        RECT 230.790 81.520 231.960 81.690 ;
        RECT 230.790 81.480 231.120 81.520 ;
        RECT 231.230 81.260 231.460 81.350 ;
        RECT 229.825 81.020 231.460 81.260 ;
        RECT 231.630 81.020 231.960 81.520 ;
        RECT 225.210 79.310 225.540 79.805 ;
        RECT 225.715 79.480 225.965 79.940 ;
        RECT 226.135 79.310 226.410 79.970 ;
        RECT 226.580 79.310 226.870 80.035 ;
        RECT 227.040 79.310 228.710 80.080 ;
        RECT 228.900 79.890 229.070 81.020 ;
        RECT 232.130 80.850 232.300 81.690 ;
        RECT 229.240 80.680 232.300 80.850 ;
        RECT 229.240 80.130 229.410 80.680 ;
        RECT 229.640 80.300 230.005 80.500 ;
        RECT 230.175 80.300 230.505 80.500 ;
        RECT 229.240 79.960 230.040 80.130 ;
        RECT 228.900 79.820 229.085 79.890 ;
        RECT 228.900 79.810 229.110 79.820 ;
        RECT 228.900 79.480 229.155 79.810 ;
        RECT 229.370 79.310 229.700 79.790 ;
        RECT 229.870 79.730 230.040 79.960 ;
        RECT 230.220 79.900 230.505 80.300 ;
        RECT 230.775 80.300 231.250 80.500 ;
        RECT 231.420 80.300 231.865 80.500 ;
        RECT 232.035 80.300 232.385 80.510 ;
        RECT 230.775 79.900 231.055 80.300 ;
        RECT 231.235 79.960 232.300 80.130 ;
        RECT 231.235 79.730 231.405 79.960 ;
        RECT 229.870 79.480 231.405 79.730 ;
        RECT 231.630 79.310 231.960 79.790 ;
        RECT 232.130 79.480 232.300 79.960 ;
        RECT 232.570 79.490 232.830 81.680 ;
        RECT 233.000 81.130 233.340 81.860 ;
        RECT 233.520 80.950 233.790 81.680 ;
        RECT 233.020 80.730 233.790 80.950 ;
        RECT 233.970 80.970 234.200 81.680 ;
        RECT 234.370 81.150 234.700 81.860 ;
        RECT 234.870 80.970 235.130 81.680 ;
        RECT 233.970 80.730 235.130 80.970 ;
        RECT 235.320 80.770 238.830 81.860 ;
        RECT 233.020 80.060 233.310 80.730 ;
        RECT 233.490 80.240 233.955 80.550 ;
        RECT 234.135 80.240 234.660 80.550 ;
        RECT 233.020 79.860 234.250 80.060 ;
        RECT 233.090 79.310 233.760 79.680 ;
        RECT 233.940 79.490 234.250 79.860 ;
        RECT 234.430 79.600 234.660 80.240 ;
        RECT 234.840 80.220 235.140 80.550 ;
        RECT 235.320 80.080 236.970 80.600 ;
        RECT 237.140 80.250 238.830 80.770 ;
        RECT 239.465 81.470 239.800 81.690 ;
        RECT 240.805 81.480 241.160 81.860 ;
        RECT 239.465 80.850 239.720 81.470 ;
        RECT 239.970 81.310 240.200 81.350 ;
        RECT 241.330 81.310 241.580 81.690 ;
        RECT 239.970 81.110 241.580 81.310 ;
        RECT 239.970 81.020 240.155 81.110 ;
        RECT 240.745 81.100 241.580 81.110 ;
        RECT 241.830 81.080 242.080 81.860 ;
        RECT 242.250 81.010 242.510 81.690 ;
        RECT 240.310 80.910 240.640 80.940 ;
        RECT 240.310 80.850 242.110 80.910 ;
        RECT 239.465 80.740 242.170 80.850 ;
        RECT 239.465 80.680 240.640 80.740 ;
        RECT 241.970 80.705 242.170 80.740 ;
        RECT 239.460 80.300 239.950 80.500 ;
        RECT 240.140 80.300 240.615 80.510 ;
        RECT 234.840 79.310 235.130 80.040 ;
        RECT 235.320 79.310 238.830 80.080 ;
        RECT 239.465 79.310 239.920 80.075 ;
        RECT 240.395 79.900 240.615 80.300 ;
        RECT 240.860 80.300 241.190 80.510 ;
        RECT 240.860 79.900 241.070 80.300 ;
        RECT 241.360 80.265 241.770 80.570 ;
        RECT 242.000 80.130 242.170 80.705 ;
        RECT 241.900 80.010 242.170 80.130 ;
        RECT 241.325 79.965 242.170 80.010 ;
        RECT 241.325 79.840 242.080 79.965 ;
        RECT 241.325 79.690 241.495 79.840 ;
        RECT 242.340 79.820 242.510 81.010 ;
        RECT 242.770 80.850 242.940 81.690 ;
        RECT 243.110 81.520 244.280 81.690 ;
        RECT 243.110 81.020 243.440 81.520 ;
        RECT 243.950 81.480 244.280 81.520 ;
        RECT 244.470 81.440 244.825 81.860 ;
        RECT 243.610 81.260 243.840 81.350 ;
        RECT 244.995 81.260 245.245 81.690 ;
        RECT 243.610 81.020 245.245 81.260 ;
        RECT 245.415 81.100 245.745 81.860 ;
        RECT 245.915 81.020 246.170 81.690 ;
        RECT 242.770 80.680 245.830 80.850 ;
        RECT 242.685 80.300 243.035 80.510 ;
        RECT 243.205 80.300 243.650 80.500 ;
        RECT 243.820 80.300 244.295 80.500 ;
        RECT 242.280 79.810 242.510 79.820 ;
        RECT 240.195 79.480 241.495 79.690 ;
        RECT 241.750 79.310 242.080 79.670 ;
        RECT 242.250 79.480 242.510 79.810 ;
        RECT 242.770 79.960 243.835 80.130 ;
        RECT 242.770 79.480 242.940 79.960 ;
        RECT 243.110 79.310 243.440 79.790 ;
        RECT 243.665 79.730 243.835 79.960 ;
        RECT 244.015 79.900 244.295 80.300 ;
        RECT 244.565 80.300 244.895 80.500 ;
        RECT 245.065 80.330 245.440 80.500 ;
        RECT 245.065 80.300 245.430 80.330 ;
        RECT 244.565 79.900 244.850 80.300 ;
        RECT 245.660 80.130 245.830 80.680 ;
        RECT 245.030 79.960 245.830 80.130 ;
        RECT 245.030 79.730 245.200 79.960 ;
        RECT 246.000 79.890 246.170 81.020 ;
        RECT 246.360 80.850 246.625 81.860 ;
        RECT 246.795 81.020 247.080 81.690 ;
        RECT 246.795 80.670 246.965 81.020 ;
        RECT 247.280 81.015 247.495 81.860 ;
        RECT 247.665 81.350 248.140 81.690 ;
        RECT 248.310 81.355 248.925 81.860 ;
        RECT 248.310 81.180 248.500 81.355 ;
        RECT 247.755 80.820 247.945 81.115 ;
        RECT 248.170 80.990 248.500 81.180 ;
        RECT 248.670 80.820 248.905 81.185 ;
        RECT 246.360 80.150 246.965 80.670 ;
        RECT 247.135 80.650 248.905 80.820 ;
        RECT 247.135 80.220 247.365 80.650 ;
        RECT 245.985 79.820 246.170 79.890 ;
        RECT 245.960 79.810 246.170 79.820 ;
        RECT 243.665 79.480 245.200 79.730 ;
        RECT 245.370 79.310 245.700 79.790 ;
        RECT 245.915 79.480 246.170 79.810 ;
        RECT 246.360 79.310 246.625 79.970 ;
        RECT 246.795 79.940 246.965 80.150 ;
        RECT 247.535 79.990 247.945 80.470 ;
        RECT 246.795 79.480 247.040 79.940 ;
        RECT 247.215 79.310 247.545 79.805 ;
        RECT 247.735 79.530 247.945 79.990 ;
        RECT 248.115 79.795 248.370 80.650 ;
        RECT 249.100 80.470 249.375 81.130 ;
        RECT 249.555 80.800 249.870 81.860 ;
        RECT 250.040 80.770 251.710 81.860 ;
        RECT 248.540 80.240 249.375 80.470 ;
        RECT 248.115 79.530 248.900 79.795 ;
        RECT 249.100 79.530 249.375 80.240 ;
        RECT 249.545 79.970 249.810 80.550 ;
        RECT 250.040 80.080 250.790 80.600 ;
        RECT 250.960 80.250 251.710 80.770 ;
        RECT 252.340 80.695 252.630 81.860 ;
        RECT 252.800 80.770 254.010 81.860 ;
        RECT 249.600 79.310 249.870 79.800 ;
        RECT 250.040 79.310 251.710 80.080 ;
        RECT 252.800 80.060 253.320 80.600 ;
        RECT 253.490 80.230 254.010 80.770 ;
        RECT 254.185 81.470 254.520 81.690 ;
        RECT 255.525 81.480 255.880 81.860 ;
        RECT 254.185 80.850 254.440 81.470 ;
        RECT 254.690 81.310 254.920 81.350 ;
        RECT 256.050 81.310 256.300 81.690 ;
        RECT 254.690 81.110 256.300 81.310 ;
        RECT 254.690 81.020 254.875 81.110 ;
        RECT 255.465 81.100 256.300 81.110 ;
        RECT 256.550 81.080 256.800 81.860 ;
        RECT 256.970 81.010 257.230 81.690 ;
        RECT 255.030 80.910 255.360 80.940 ;
        RECT 255.030 80.850 256.830 80.910 ;
        RECT 254.185 80.740 256.890 80.850 ;
        RECT 254.185 80.680 255.360 80.740 ;
        RECT 256.690 80.705 256.890 80.740 ;
        RECT 254.180 80.300 254.670 80.500 ;
        RECT 254.860 80.300 255.335 80.510 ;
        RECT 252.340 79.310 252.630 80.035 ;
        RECT 252.800 79.310 254.010 80.060 ;
        RECT 254.185 79.310 254.640 80.075 ;
        RECT 255.115 79.900 255.335 80.300 ;
        RECT 255.580 80.300 255.910 80.510 ;
        RECT 255.580 79.900 255.790 80.300 ;
        RECT 256.080 80.265 256.490 80.570 ;
        RECT 256.720 80.130 256.890 80.705 ;
        RECT 256.620 80.010 256.890 80.130 ;
        RECT 256.045 79.965 256.890 80.010 ;
        RECT 256.045 79.840 256.800 79.965 ;
        RECT 256.045 79.690 256.215 79.840 ;
        RECT 257.060 79.810 257.230 81.010 ;
        RECT 257.490 80.850 257.660 81.690 ;
        RECT 257.830 81.520 259.000 81.690 ;
        RECT 257.830 81.020 258.160 81.520 ;
        RECT 258.670 81.480 259.000 81.520 ;
        RECT 259.190 81.440 259.545 81.860 ;
        RECT 258.330 81.260 258.560 81.350 ;
        RECT 259.715 81.260 259.965 81.690 ;
        RECT 258.330 81.020 259.965 81.260 ;
        RECT 260.135 81.100 260.465 81.860 ;
        RECT 260.635 81.020 260.890 81.690 ;
        RECT 257.490 80.680 260.550 80.850 ;
        RECT 257.405 80.300 257.755 80.510 ;
        RECT 257.925 80.300 258.370 80.500 ;
        RECT 258.540 80.300 259.015 80.500 ;
        RECT 254.915 79.480 256.215 79.690 ;
        RECT 256.470 79.310 256.800 79.670 ;
        RECT 256.970 79.480 257.230 79.810 ;
        RECT 257.490 79.960 258.555 80.130 ;
        RECT 257.490 79.480 257.660 79.960 ;
        RECT 257.830 79.310 258.160 79.790 ;
        RECT 258.385 79.730 258.555 79.960 ;
        RECT 258.735 79.900 259.015 80.300 ;
        RECT 259.285 80.300 259.615 80.500 ;
        RECT 259.785 80.300 260.150 80.500 ;
        RECT 259.285 79.900 259.570 80.300 ;
        RECT 260.380 80.130 260.550 80.680 ;
        RECT 259.750 79.960 260.550 80.130 ;
        RECT 259.750 79.730 259.920 79.960 ;
        RECT 260.720 79.890 260.890 81.020 ;
        RECT 260.705 79.820 260.890 79.890 ;
        RECT 260.680 79.810 260.890 79.820 ;
        RECT 258.385 79.480 259.920 79.730 ;
        RECT 260.090 79.310 260.420 79.790 ;
        RECT 260.635 79.480 260.890 79.810 ;
        RECT 261.100 81.020 261.355 81.690 ;
        RECT 261.525 81.100 261.855 81.860 ;
        RECT 262.025 81.260 262.275 81.690 ;
        RECT 262.445 81.440 262.800 81.860 ;
        RECT 262.990 81.520 264.160 81.690 ;
        RECT 262.990 81.480 263.320 81.520 ;
        RECT 263.430 81.260 263.660 81.350 ;
        RECT 262.025 81.020 263.660 81.260 ;
        RECT 263.830 81.020 264.160 81.520 ;
        RECT 261.100 81.010 261.310 81.020 ;
        RECT 261.100 79.890 261.270 81.010 ;
        RECT 264.330 80.850 264.500 81.690 ;
        RECT 261.440 80.680 264.500 80.850 ;
        RECT 264.760 81.010 265.020 81.690 ;
        RECT 265.190 81.080 265.440 81.860 ;
        RECT 265.690 81.310 265.940 81.690 ;
        RECT 266.110 81.480 266.465 81.860 ;
        RECT 267.470 81.470 267.805 81.690 ;
        RECT 267.070 81.310 267.300 81.350 ;
        RECT 265.690 81.110 267.300 81.310 ;
        RECT 265.690 81.100 266.525 81.110 ;
        RECT 267.115 81.020 267.300 81.110 ;
        RECT 261.440 80.130 261.610 80.680 ;
        RECT 261.830 80.330 262.205 80.500 ;
        RECT 261.840 80.300 262.205 80.330 ;
        RECT 262.375 80.300 262.705 80.500 ;
        RECT 261.440 79.960 262.240 80.130 ;
        RECT 261.100 79.810 261.285 79.890 ;
        RECT 261.100 79.480 261.355 79.810 ;
        RECT 261.570 79.310 261.900 79.790 ;
        RECT 262.070 79.730 262.240 79.960 ;
        RECT 262.420 79.900 262.705 80.300 ;
        RECT 262.975 80.300 263.450 80.500 ;
        RECT 263.620 80.300 264.065 80.500 ;
        RECT 264.235 80.300 264.585 80.510 ;
        RECT 262.975 79.900 263.255 80.300 ;
        RECT 263.435 79.960 264.500 80.130 ;
        RECT 263.435 79.730 263.605 79.960 ;
        RECT 262.070 79.480 263.605 79.730 ;
        RECT 263.830 79.310 264.160 79.790 ;
        RECT 264.330 79.480 264.500 79.960 ;
        RECT 264.760 79.810 264.930 81.010 ;
        RECT 266.630 80.910 266.960 80.940 ;
        RECT 265.160 80.850 266.960 80.910 ;
        RECT 267.550 80.850 267.805 81.470 ;
        RECT 267.985 81.350 269.640 81.640 ;
        RECT 265.100 80.740 267.805 80.850 ;
        RECT 265.100 80.705 265.300 80.740 ;
        RECT 265.100 80.130 265.270 80.705 ;
        RECT 266.630 80.680 267.805 80.740 ;
        RECT 267.985 81.010 269.575 81.180 ;
        RECT 269.810 81.060 270.090 81.860 ;
        RECT 267.985 80.720 268.305 81.010 ;
        RECT 269.405 80.890 269.575 81.010 ;
        RECT 268.500 80.670 269.215 80.840 ;
        RECT 269.405 80.720 270.130 80.890 ;
        RECT 270.300 80.720 270.570 81.690 ;
        RECT 270.740 81.425 276.085 81.860 ;
        RECT 265.500 80.265 265.910 80.570 ;
        RECT 266.080 80.300 266.410 80.510 ;
        RECT 265.100 80.010 265.370 80.130 ;
        RECT 265.100 79.965 265.945 80.010 ;
        RECT 265.190 79.840 265.945 79.965 ;
        RECT 266.200 79.900 266.410 80.300 ;
        RECT 266.655 80.300 267.130 80.510 ;
        RECT 267.320 80.300 267.810 80.500 ;
        RECT 266.655 79.900 266.875 80.300 ;
        RECT 264.760 79.480 265.020 79.810 ;
        RECT 265.775 79.690 265.945 79.840 ;
        RECT 265.190 79.310 265.520 79.670 ;
        RECT 265.775 79.480 267.075 79.690 ;
        RECT 267.350 79.310 267.805 80.075 ;
        RECT 267.985 79.980 268.335 80.550 ;
        RECT 268.505 80.220 269.215 80.670 ;
        RECT 269.960 80.550 270.130 80.720 ;
        RECT 269.385 80.220 269.790 80.550 ;
        RECT 269.960 80.220 270.230 80.550 ;
        RECT 269.960 80.050 270.130 80.220 ;
        RECT 268.520 79.880 270.130 80.050 ;
        RECT 270.400 79.985 270.570 80.720 ;
        RECT 267.990 79.310 268.320 79.810 ;
        RECT 268.520 79.530 268.690 79.880 ;
        RECT 268.890 79.310 269.220 79.710 ;
        RECT 269.390 79.530 269.560 79.880 ;
        RECT 269.730 79.310 270.110 79.710 ;
        RECT 270.300 79.640 270.570 79.985 ;
        RECT 272.325 79.855 272.665 80.685 ;
        RECT 274.145 80.175 274.495 81.425 ;
        RECT 276.260 80.770 277.930 81.860 ;
        RECT 276.260 80.080 277.010 80.600 ;
        RECT 277.180 80.250 277.930 80.770 ;
        RECT 278.100 80.695 278.390 81.860 ;
        RECT 278.560 80.770 280.230 81.860 ;
        RECT 278.560 80.080 279.310 80.600 ;
        RECT 279.480 80.250 280.230 80.770 ;
        RECT 280.865 80.720 281.200 81.690 ;
        RECT 281.370 80.720 281.540 81.860 ;
        RECT 281.710 81.520 283.740 81.690 ;
        RECT 270.740 79.310 276.085 79.855 ;
        RECT 276.260 79.310 277.930 80.080 ;
        RECT 278.100 79.310 278.390 80.035 ;
        RECT 278.560 79.310 280.230 80.080 ;
        RECT 280.865 80.050 281.035 80.720 ;
        RECT 281.710 80.550 281.880 81.520 ;
        RECT 281.205 80.220 281.460 80.550 ;
        RECT 281.685 80.220 281.880 80.550 ;
        RECT 282.050 81.180 283.175 81.350 ;
        RECT 281.290 80.050 281.460 80.220 ;
        RECT 282.050 80.050 282.220 81.180 ;
        RECT 280.865 79.480 281.120 80.050 ;
        RECT 281.290 79.880 282.220 80.050 ;
        RECT 282.390 80.840 283.400 81.010 ;
        RECT 282.390 80.040 282.560 80.840 ;
        RECT 282.045 79.845 282.220 79.880 ;
        RECT 281.290 79.310 281.620 79.710 ;
        RECT 282.045 79.480 282.575 79.845 ;
        RECT 282.765 79.820 283.040 80.640 ;
        RECT 282.760 79.650 283.040 79.820 ;
        RECT 282.765 79.480 283.040 79.650 ;
        RECT 283.210 79.480 283.400 80.840 ;
        RECT 283.570 80.855 283.740 81.520 ;
        RECT 283.910 81.100 284.080 81.860 ;
        RECT 284.315 81.100 284.830 81.510 ;
        RECT 283.570 80.665 284.320 80.855 ;
        RECT 284.490 80.290 284.830 81.100 ;
        RECT 283.600 80.120 284.830 80.290 ;
        RECT 285.005 80.720 285.340 81.690 ;
        RECT 285.510 80.720 285.680 81.860 ;
        RECT 285.850 81.520 287.880 81.690 ;
        RECT 283.580 79.310 284.090 79.845 ;
        RECT 284.310 79.515 284.555 80.120 ;
        RECT 285.005 80.050 285.175 80.720 ;
        RECT 285.850 80.550 286.020 81.520 ;
        RECT 285.345 80.220 285.600 80.550 ;
        RECT 285.825 80.220 286.020 80.550 ;
        RECT 286.190 81.180 287.315 81.350 ;
        RECT 285.430 80.050 285.600 80.220 ;
        RECT 286.190 80.050 286.360 81.180 ;
        RECT 285.005 79.480 285.260 80.050 ;
        RECT 285.430 79.880 286.360 80.050 ;
        RECT 286.530 80.840 287.540 81.010 ;
        RECT 286.530 80.040 286.700 80.840 ;
        RECT 286.185 79.845 286.360 79.880 ;
        RECT 285.430 79.310 285.760 79.710 ;
        RECT 286.185 79.480 286.715 79.845 ;
        RECT 286.905 79.820 287.180 80.640 ;
        RECT 286.900 79.650 287.180 79.820 ;
        RECT 286.905 79.480 287.180 79.650 ;
        RECT 287.350 79.480 287.540 80.840 ;
        RECT 287.710 80.855 287.880 81.520 ;
        RECT 288.050 81.100 288.220 81.860 ;
        RECT 288.455 81.100 288.970 81.510 ;
        RECT 287.710 80.665 288.460 80.855 ;
        RECT 288.630 80.290 288.970 81.100 ;
        RECT 289.140 80.770 290.350 81.860 ;
        RECT 287.740 80.120 288.970 80.290 ;
        RECT 287.720 79.310 288.230 79.845 ;
        RECT 288.450 79.515 288.695 80.120 ;
        RECT 289.140 80.060 289.660 80.600 ;
        RECT 289.830 80.230 290.350 80.770 ;
        RECT 290.520 81.100 291.035 81.510 ;
        RECT 291.270 81.100 291.440 81.860 ;
        RECT 291.610 81.520 293.640 81.690 ;
        RECT 290.520 80.290 290.860 81.100 ;
        RECT 291.610 80.855 291.780 81.520 ;
        RECT 292.175 81.180 293.300 81.350 ;
        RECT 291.030 80.665 291.780 80.855 ;
        RECT 291.950 80.840 292.960 81.010 ;
        RECT 290.520 80.120 291.750 80.290 ;
        RECT 289.140 79.310 290.350 80.060 ;
        RECT 290.795 79.515 291.040 80.120 ;
        RECT 291.260 79.310 291.770 79.845 ;
        RECT 291.950 79.480 292.140 80.840 ;
        RECT 292.310 79.820 292.585 80.640 ;
        RECT 292.790 80.040 292.960 80.840 ;
        RECT 293.130 80.050 293.300 81.180 ;
        RECT 293.470 80.550 293.640 81.520 ;
        RECT 293.810 80.720 293.980 81.860 ;
        RECT 294.150 80.720 294.485 81.690 ;
        RECT 293.470 80.220 293.665 80.550 ;
        RECT 293.890 80.220 294.145 80.550 ;
        RECT 293.890 80.050 294.060 80.220 ;
        RECT 294.315 80.050 294.485 80.720 ;
        RECT 293.130 79.880 294.060 80.050 ;
        RECT 293.130 79.845 293.305 79.880 ;
        RECT 292.310 79.650 292.590 79.820 ;
        RECT 292.310 79.480 292.585 79.650 ;
        RECT 292.775 79.480 293.305 79.845 ;
        RECT 293.730 79.310 294.060 79.710 ;
        RECT 294.230 79.480 294.485 80.050 ;
        RECT 294.665 80.670 294.920 81.550 ;
        RECT 295.090 80.720 295.395 81.860 ;
        RECT 295.735 81.480 296.065 81.860 ;
        RECT 296.245 81.310 296.415 81.600 ;
        RECT 296.585 81.400 296.835 81.860 ;
        RECT 295.615 81.140 296.415 81.310 ;
        RECT 297.005 81.350 297.875 81.690 ;
        RECT 294.665 80.020 294.875 80.670 ;
        RECT 295.615 80.550 295.785 81.140 ;
        RECT 297.005 80.970 297.175 81.350 ;
        RECT 298.110 81.230 298.280 81.690 ;
        RECT 298.450 81.400 298.820 81.860 ;
        RECT 299.115 81.260 299.285 81.600 ;
        RECT 299.455 81.430 299.785 81.860 ;
        RECT 300.020 81.260 300.190 81.600 ;
        RECT 295.955 80.800 297.175 80.970 ;
        RECT 297.345 80.890 297.805 81.180 ;
        RECT 298.110 81.060 298.670 81.230 ;
        RECT 299.115 81.090 300.190 81.260 ;
        RECT 300.360 81.360 301.040 81.690 ;
        RECT 301.255 81.360 301.505 81.690 ;
        RECT 301.675 81.400 301.925 81.860 ;
        RECT 298.500 80.920 298.670 81.060 ;
        RECT 297.345 80.880 298.310 80.890 ;
        RECT 297.005 80.710 297.175 80.800 ;
        RECT 297.635 80.720 298.310 80.880 ;
        RECT 295.045 80.520 295.785 80.550 ;
        RECT 295.045 80.220 295.960 80.520 ;
        RECT 295.635 80.045 295.960 80.220 ;
        RECT 294.665 79.490 294.920 80.020 ;
        RECT 295.090 79.310 295.395 79.770 ;
        RECT 295.640 79.690 295.960 80.045 ;
        RECT 296.130 80.260 296.670 80.630 ;
        RECT 297.005 80.540 297.410 80.710 ;
        RECT 296.130 79.860 296.370 80.260 ;
        RECT 296.850 80.090 297.070 80.370 ;
        RECT 296.540 79.920 297.070 80.090 ;
        RECT 296.540 79.690 296.710 79.920 ;
        RECT 297.240 79.760 297.410 80.540 ;
        RECT 297.580 79.930 297.930 80.550 ;
        RECT 298.100 79.930 298.310 80.720 ;
        RECT 298.500 80.750 300.000 80.920 ;
        RECT 298.500 80.060 298.670 80.750 ;
        RECT 300.360 80.580 300.530 81.360 ;
        RECT 301.335 81.230 301.505 81.360 ;
        RECT 298.840 80.410 300.530 80.580 ;
        RECT 300.700 80.800 301.165 81.190 ;
        RECT 301.335 81.060 301.730 81.230 ;
        RECT 298.840 80.230 299.010 80.410 ;
        RECT 295.640 79.520 296.710 79.690 ;
        RECT 296.880 79.310 297.070 79.750 ;
        RECT 297.240 79.480 298.190 79.760 ;
        RECT 298.500 79.670 298.760 80.060 ;
        RECT 299.180 79.990 299.970 80.240 ;
        RECT 298.410 79.500 298.760 79.670 ;
        RECT 298.970 79.310 299.300 79.770 ;
        RECT 300.175 79.700 300.345 80.410 ;
        RECT 300.700 80.210 300.870 80.800 ;
        RECT 300.515 79.990 300.870 80.210 ;
        RECT 301.040 79.990 301.390 80.610 ;
        RECT 301.560 79.700 301.730 81.060 ;
        RECT 302.095 80.890 302.420 81.675 ;
        RECT 301.900 79.840 302.360 80.890 ;
        RECT 300.175 79.530 301.030 79.700 ;
        RECT 301.235 79.530 301.730 79.700 ;
        RECT 301.900 79.310 302.230 79.670 ;
        RECT 302.590 79.570 302.760 81.690 ;
        RECT 302.930 81.360 303.260 81.860 ;
        RECT 303.430 81.190 303.685 81.690 ;
        RECT 302.935 81.020 303.685 81.190 ;
        RECT 302.935 80.030 303.165 81.020 ;
        RECT 303.335 80.200 303.685 80.850 ;
        RECT 303.860 80.695 304.150 81.860 ;
        RECT 304.320 81.425 309.665 81.860 ;
        RECT 302.935 79.860 303.685 80.030 ;
        RECT 302.930 79.310 303.260 79.690 ;
        RECT 303.430 79.570 303.685 79.860 ;
        RECT 303.860 79.310 304.150 80.035 ;
        RECT 305.905 79.855 306.245 80.685 ;
        RECT 307.725 80.175 308.075 81.425 ;
        RECT 309.840 80.770 311.050 81.860 ;
        RECT 309.840 80.230 310.360 80.770 ;
        RECT 310.530 80.060 311.050 80.600 ;
        RECT 304.320 79.310 309.665 79.855 ;
        RECT 309.840 79.310 311.050 80.060 ;
        RECT 162.095 79.140 311.135 79.310 ;
        RECT 162.180 78.390 163.390 79.140 ;
        RECT 163.560 78.595 168.905 79.140 ;
        RECT 162.180 77.850 162.700 78.390 ;
        RECT 162.870 77.680 163.390 78.220 ;
        RECT 165.145 77.765 165.485 78.595 ;
        RECT 170.005 78.590 170.260 78.880 ;
        RECT 170.430 78.760 170.760 79.140 ;
        RECT 170.005 78.420 170.755 78.590 ;
        RECT 162.180 76.590 163.390 77.680 ;
        RECT 166.965 77.025 167.315 78.275 ;
        RECT 170.005 77.600 170.355 78.250 ;
        RECT 170.525 77.430 170.755 78.420 ;
        RECT 170.005 77.260 170.755 77.430 ;
        RECT 163.560 76.590 168.905 77.025 ;
        RECT 170.005 76.760 170.260 77.260 ;
        RECT 170.430 76.590 170.760 77.090 ;
        RECT 170.930 76.760 171.100 78.880 ;
        RECT 171.460 78.780 171.790 79.140 ;
        RECT 171.960 78.750 172.455 78.920 ;
        RECT 172.660 78.750 173.515 78.920 ;
        RECT 171.330 77.560 171.790 78.610 ;
        RECT 171.270 76.775 171.595 77.560 ;
        RECT 171.960 77.390 172.130 78.750 ;
        RECT 172.300 77.840 172.650 78.460 ;
        RECT 172.820 78.240 173.175 78.460 ;
        RECT 172.820 77.650 172.990 78.240 ;
        RECT 173.345 78.040 173.515 78.750 ;
        RECT 174.390 78.680 174.720 79.140 ;
        RECT 174.930 78.780 175.280 78.950 ;
        RECT 173.720 78.210 174.510 78.460 ;
        RECT 174.930 78.390 175.190 78.780 ;
        RECT 175.500 78.690 176.450 78.970 ;
        RECT 176.620 78.700 176.810 79.140 ;
        RECT 176.980 78.760 178.050 78.930 ;
        RECT 174.680 78.040 174.850 78.220 ;
        RECT 171.960 77.220 172.355 77.390 ;
        RECT 172.525 77.260 172.990 77.650 ;
        RECT 173.160 77.870 174.850 78.040 ;
        RECT 172.185 77.090 172.355 77.220 ;
        RECT 173.160 77.090 173.330 77.870 ;
        RECT 175.020 77.700 175.190 78.390 ;
        RECT 173.690 77.530 175.190 77.700 ;
        RECT 175.380 77.730 175.590 78.520 ;
        RECT 175.760 77.900 176.110 78.520 ;
        RECT 176.280 77.910 176.450 78.690 ;
        RECT 176.980 78.530 177.150 78.760 ;
        RECT 176.620 78.360 177.150 78.530 ;
        RECT 176.620 78.080 176.840 78.360 ;
        RECT 177.320 78.190 177.560 78.590 ;
        RECT 176.280 77.740 176.685 77.910 ;
        RECT 177.020 77.820 177.560 78.190 ;
        RECT 177.730 78.405 178.050 78.760 ;
        RECT 178.295 78.680 178.600 79.140 ;
        RECT 178.770 78.430 179.020 78.960 ;
        RECT 177.730 78.230 178.055 78.405 ;
        RECT 177.730 77.930 178.645 78.230 ;
        RECT 177.905 77.900 178.645 77.930 ;
        RECT 175.380 77.570 176.055 77.730 ;
        RECT 176.515 77.650 176.685 77.740 ;
        RECT 175.380 77.560 176.345 77.570 ;
        RECT 175.020 77.390 175.190 77.530 ;
        RECT 171.765 76.590 172.015 77.050 ;
        RECT 172.185 76.760 172.435 77.090 ;
        RECT 172.650 76.760 173.330 77.090 ;
        RECT 173.500 77.190 174.575 77.360 ;
        RECT 175.020 77.220 175.580 77.390 ;
        RECT 175.885 77.270 176.345 77.560 ;
        RECT 176.515 77.480 177.735 77.650 ;
        RECT 173.500 76.850 173.670 77.190 ;
        RECT 173.905 76.590 174.235 77.020 ;
        RECT 174.405 76.850 174.575 77.190 ;
        RECT 174.870 76.590 175.240 77.050 ;
        RECT 175.410 76.760 175.580 77.220 ;
        RECT 176.515 77.100 176.685 77.480 ;
        RECT 177.905 77.310 178.075 77.900 ;
        RECT 178.815 77.780 179.020 78.430 ;
        RECT 179.190 78.385 179.440 79.140 ;
        RECT 179.665 78.400 179.920 78.970 ;
        RECT 180.090 78.740 180.420 79.140 ;
        RECT 180.845 78.605 181.375 78.970 ;
        RECT 180.845 78.570 181.020 78.605 ;
        RECT 180.090 78.400 181.020 78.570 ;
        RECT 175.815 76.760 176.685 77.100 ;
        RECT 177.275 77.140 178.075 77.310 ;
        RECT 176.855 76.590 177.105 77.050 ;
        RECT 177.275 76.850 177.445 77.140 ;
        RECT 177.625 76.590 177.955 76.970 ;
        RECT 178.295 76.590 178.600 77.730 ;
        RECT 178.770 76.900 179.020 77.780 ;
        RECT 179.665 77.730 179.835 78.400 ;
        RECT 180.090 78.230 180.260 78.400 ;
        RECT 180.005 77.900 180.260 78.230 ;
        RECT 180.485 77.900 180.680 78.230 ;
        RECT 179.190 76.590 179.440 77.730 ;
        RECT 179.665 76.760 180.000 77.730 ;
        RECT 180.170 76.590 180.340 77.730 ;
        RECT 180.510 76.930 180.680 77.900 ;
        RECT 180.850 77.270 181.020 78.400 ;
        RECT 181.190 77.610 181.360 78.410 ;
        RECT 181.565 78.120 181.840 78.970 ;
        RECT 181.560 77.950 181.840 78.120 ;
        RECT 181.565 77.810 181.840 77.950 ;
        RECT 182.010 77.610 182.200 78.970 ;
        RECT 182.380 78.605 182.890 79.140 ;
        RECT 183.110 78.330 183.355 78.935 ;
        RECT 184.740 78.510 185.070 78.970 ;
        RECT 185.250 78.680 185.420 79.140 ;
        RECT 185.600 78.510 185.930 78.970 ;
        RECT 186.160 78.680 186.330 79.140 ;
        RECT 186.570 78.800 187.760 78.970 ;
        RECT 186.570 78.510 186.900 78.800 ;
        RECT 187.450 78.630 187.760 78.800 ;
        RECT 184.740 78.340 186.900 78.510 ;
        RECT 182.400 78.160 183.630 78.330 ;
        RECT 181.190 77.440 182.200 77.610 ;
        RECT 182.370 77.595 183.120 77.785 ;
        RECT 180.850 77.100 181.975 77.270 ;
        RECT 182.370 76.930 182.540 77.595 ;
        RECT 183.290 77.350 183.630 78.160 ;
        RECT 184.755 77.780 185.085 78.170 ;
        RECT 185.255 77.950 186.055 78.150 ;
        RECT 186.235 77.780 186.730 78.150 ;
        RECT 184.755 77.610 186.730 77.780 ;
        RECT 187.070 77.440 187.280 78.630 ;
        RECT 187.450 77.825 187.765 78.460 ;
        RECT 187.940 78.415 188.230 79.140 ;
        RECT 189.105 78.660 189.405 79.140 ;
        RECT 189.575 78.490 189.835 78.945 ;
        RECT 190.005 78.660 190.265 79.140 ;
        RECT 190.435 78.490 190.695 78.945 ;
        RECT 190.865 78.660 191.125 79.140 ;
        RECT 191.295 78.490 191.555 78.945 ;
        RECT 191.725 78.660 191.985 79.140 ;
        RECT 192.155 78.490 192.415 78.945 ;
        RECT 192.585 78.615 192.845 79.140 ;
        RECT 189.105 78.320 192.415 78.490 ;
        RECT 180.510 76.760 182.540 76.930 ;
        RECT 182.710 76.590 182.880 77.350 ;
        RECT 183.115 76.940 183.630 77.350 ;
        RECT 184.740 76.590 185.070 77.440 ;
        RECT 185.240 76.930 185.460 77.440 ;
        RECT 185.630 77.260 187.280 77.440 ;
        RECT 185.630 77.100 185.930 77.260 ;
        RECT 186.160 76.930 186.350 77.090 ;
        RECT 185.240 76.760 186.350 76.930 ;
        RECT 186.545 76.590 186.875 77.050 ;
        RECT 187.045 76.760 187.280 77.260 ;
        RECT 187.450 76.590 187.760 77.655 ;
        RECT 187.940 76.590 188.230 77.755 ;
        RECT 189.105 77.730 190.075 78.320 ;
        RECT 193.015 78.150 193.265 78.960 ;
        RECT 193.445 78.680 193.690 79.140 ;
        RECT 193.940 78.570 194.195 78.920 ;
        RECT 194.365 78.740 194.695 79.140 ;
        RECT 194.865 78.570 195.035 78.920 ;
        RECT 195.205 78.740 195.585 79.140 ;
        RECT 190.245 77.900 193.265 78.150 ;
        RECT 193.435 77.900 193.750 78.510 ;
        RECT 193.940 78.400 195.605 78.570 ;
        RECT 195.775 78.465 196.050 78.810 ;
        RECT 195.435 78.230 195.605 78.400 ;
        RECT 193.920 77.900 194.270 78.230 ;
        RECT 194.440 77.900 195.265 78.230 ;
        RECT 195.435 77.900 195.710 78.230 ;
        RECT 189.105 77.490 192.415 77.730 ;
        RECT 189.110 76.590 189.405 77.320 ;
        RECT 189.575 76.765 189.835 77.490 ;
        RECT 190.005 76.590 190.265 77.320 ;
        RECT 190.435 76.765 190.695 77.490 ;
        RECT 190.865 76.590 191.125 77.320 ;
        RECT 191.295 76.765 191.555 77.490 ;
        RECT 191.725 76.590 191.985 77.320 ;
        RECT 192.155 76.765 192.415 77.490 ;
        RECT 192.585 76.590 192.845 77.700 ;
        RECT 193.015 76.765 193.265 77.900 ;
        RECT 193.445 76.590 193.740 77.700 ;
        RECT 193.940 77.440 194.270 77.730 ;
        RECT 194.440 77.610 194.665 77.900 ;
        RECT 195.435 77.730 195.605 77.900 ;
        RECT 195.880 77.730 196.050 78.465 ;
        RECT 196.220 78.310 196.510 79.140 ;
        RECT 196.885 78.360 197.385 78.970 ;
        RECT 196.680 77.900 197.030 78.150 ;
        RECT 194.935 77.560 195.605 77.730 ;
        RECT 194.935 77.440 195.105 77.560 ;
        RECT 193.940 77.270 195.105 77.440 ;
        RECT 193.920 76.810 195.115 77.100 ;
        RECT 195.285 76.590 195.565 77.390 ;
        RECT 195.775 76.760 196.050 77.730 ;
        RECT 196.220 76.590 196.510 77.795 ;
        RECT 197.215 77.730 197.385 78.360 ;
        RECT 198.015 78.490 198.345 78.970 ;
        RECT 198.515 78.680 198.740 79.140 ;
        RECT 198.910 78.490 199.240 78.970 ;
        RECT 198.015 78.320 199.240 78.490 ;
        RECT 199.430 78.340 199.680 79.140 ;
        RECT 199.850 78.340 200.190 78.970 ;
        RECT 197.555 77.950 197.885 78.150 ;
        RECT 198.055 77.950 198.385 78.150 ;
        RECT 198.555 77.950 198.975 78.150 ;
        RECT 199.150 77.980 199.845 78.150 ;
        RECT 199.150 77.730 199.320 77.980 ;
        RECT 200.015 77.730 200.190 78.340 ;
        RECT 200.360 78.370 203.870 79.140 ;
        RECT 204.500 78.650 204.770 79.140 ;
        RECT 200.360 77.850 202.010 78.370 ;
        RECT 196.885 77.560 199.320 77.730 ;
        RECT 196.885 76.760 197.215 77.560 ;
        RECT 197.385 76.590 197.715 77.390 ;
        RECT 198.015 76.760 198.345 77.560 ;
        RECT 198.990 76.590 199.240 77.390 ;
        RECT 199.510 76.590 199.680 77.730 ;
        RECT 199.850 76.760 200.190 77.730 ;
        RECT 202.180 77.680 203.870 78.200 ;
        RECT 204.560 77.900 204.825 78.480 ;
        RECT 204.995 78.210 205.270 78.920 ;
        RECT 205.470 78.655 206.255 78.920 ;
        RECT 204.995 77.980 205.830 78.210 ;
        RECT 200.360 76.590 203.870 77.680 ;
        RECT 204.500 76.590 204.815 77.650 ;
        RECT 204.995 77.320 205.270 77.980 ;
        RECT 206.000 77.800 206.255 78.655 ;
        RECT 206.425 78.460 206.635 78.920 ;
        RECT 206.825 78.645 207.155 79.140 ;
        RECT 207.330 78.510 207.575 78.970 ;
        RECT 206.425 77.980 206.835 78.460 ;
        RECT 207.405 78.300 207.575 78.510 ;
        RECT 207.745 78.480 208.010 79.140 ;
        RECT 208.180 78.370 210.770 79.140 ;
        RECT 211.105 78.630 211.345 79.140 ;
        RECT 211.525 78.630 211.805 78.960 ;
        RECT 212.035 78.630 212.250 79.140 ;
        RECT 207.005 77.800 207.235 78.230 ;
        RECT 205.465 77.630 207.235 77.800 ;
        RECT 207.405 77.780 208.010 78.300 ;
        RECT 208.180 77.850 209.390 78.370 ;
        RECT 205.465 77.265 205.700 77.630 ;
        RECT 205.870 77.270 206.200 77.460 ;
        RECT 206.425 77.335 206.615 77.630 ;
        RECT 205.870 77.095 206.060 77.270 ;
        RECT 205.445 76.590 206.060 77.095 ;
        RECT 206.230 76.760 206.705 77.100 ;
        RECT 206.875 76.590 207.090 77.435 ;
        RECT 207.405 77.430 207.575 77.780 ;
        RECT 209.560 77.680 210.770 78.200 ;
        RECT 211.000 77.900 211.355 78.460 ;
        RECT 211.525 77.730 211.695 78.630 ;
        RECT 211.865 77.900 212.130 78.460 ;
        RECT 212.420 78.400 213.035 78.970 ;
        RECT 213.700 78.415 213.990 79.140 ;
        RECT 214.160 78.595 219.505 79.140 ;
        RECT 212.380 77.730 212.550 78.230 ;
        RECT 207.290 76.760 207.575 77.430 ;
        RECT 207.745 76.590 208.010 77.600 ;
        RECT 208.180 76.590 210.770 77.680 ;
        RECT 211.125 77.560 212.550 77.730 ;
        RECT 211.125 77.385 211.515 77.560 ;
        RECT 212.000 76.590 212.330 77.390 ;
        RECT 212.720 77.380 213.035 78.400 ;
        RECT 215.745 77.765 216.085 78.595 ;
        RECT 219.680 78.370 223.190 79.140 ;
        RECT 212.500 76.760 213.035 77.380 ;
        RECT 213.700 76.590 213.990 77.755 ;
        RECT 217.565 77.025 217.915 78.275 ;
        RECT 219.680 77.850 221.330 78.370 ;
        RECT 221.500 77.680 223.190 78.200 ;
        RECT 214.160 76.590 219.505 77.025 ;
        RECT 219.680 76.590 223.190 77.680 ;
        RECT 223.820 78.195 224.160 78.970 ;
        RECT 224.330 78.680 224.500 79.140 ;
        RECT 224.740 78.705 225.100 78.970 ;
        RECT 224.740 78.700 225.095 78.705 ;
        RECT 224.740 78.690 225.090 78.700 ;
        RECT 224.740 78.685 225.085 78.690 ;
        RECT 224.740 78.675 225.080 78.685 ;
        RECT 225.730 78.680 225.900 79.140 ;
        RECT 224.740 78.670 225.075 78.675 ;
        RECT 224.740 78.660 225.065 78.670 ;
        RECT 224.740 78.650 225.055 78.660 ;
        RECT 224.740 78.510 225.040 78.650 ;
        RECT 224.330 78.320 225.040 78.510 ;
        RECT 225.230 78.510 225.560 78.590 ;
        RECT 226.070 78.510 226.410 78.970 ;
        RECT 227.040 78.650 227.310 79.140 ;
        RECT 225.230 78.320 226.410 78.510 ;
        RECT 223.820 76.760 224.100 78.195 ;
        RECT 224.330 77.750 224.615 78.320 ;
        RECT 224.800 77.920 225.270 78.150 ;
        RECT 225.440 78.130 225.770 78.150 ;
        RECT 225.440 77.950 225.890 78.130 ;
        RECT 226.080 77.950 226.410 78.150 ;
        RECT 224.330 77.535 225.480 77.750 ;
        RECT 224.270 76.590 224.980 77.365 ;
        RECT 225.150 76.760 225.480 77.535 ;
        RECT 225.675 76.835 225.890 77.950 ;
        RECT 226.180 77.610 226.410 77.950 ;
        RECT 227.100 77.900 227.365 78.480 ;
        RECT 227.535 78.210 227.810 78.920 ;
        RECT 228.010 78.655 228.795 78.920 ;
        RECT 227.535 77.980 228.370 78.210 ;
        RECT 226.070 76.590 226.400 77.310 ;
        RECT 227.040 76.590 227.355 77.650 ;
        RECT 227.535 77.320 227.810 77.980 ;
        RECT 228.540 77.800 228.795 78.655 ;
        RECT 228.965 78.460 229.175 78.920 ;
        RECT 229.365 78.645 229.695 79.140 ;
        RECT 229.870 78.510 230.115 78.970 ;
        RECT 228.965 77.980 229.375 78.460 ;
        RECT 229.945 78.300 230.115 78.510 ;
        RECT 230.285 78.480 230.550 79.140 ;
        RECT 230.720 78.595 236.065 79.140 ;
        RECT 229.545 77.800 229.775 78.230 ;
        RECT 228.005 77.630 229.775 77.800 ;
        RECT 229.945 77.780 230.550 78.300 ;
        RECT 228.005 77.265 228.240 77.630 ;
        RECT 228.410 77.270 228.740 77.460 ;
        RECT 228.965 77.335 229.155 77.630 ;
        RECT 228.410 77.095 228.600 77.270 ;
        RECT 227.985 76.590 228.600 77.095 ;
        RECT 228.770 76.760 229.245 77.100 ;
        RECT 229.415 76.590 229.630 77.435 ;
        RECT 229.945 77.430 230.115 77.780 ;
        RECT 232.305 77.765 232.645 78.595 ;
        RECT 236.240 78.370 238.830 79.140 ;
        RECT 239.460 78.415 239.750 79.140 ;
        RECT 239.920 78.370 242.510 79.140 ;
        RECT 242.685 78.375 243.140 79.140 ;
        RECT 243.415 78.760 244.715 78.970 ;
        RECT 244.970 78.780 245.300 79.140 ;
        RECT 244.545 78.610 244.715 78.760 ;
        RECT 245.470 78.640 245.730 78.970 ;
        RECT 245.910 78.640 246.240 79.140 ;
        RECT 229.830 76.760 230.115 77.430 ;
        RECT 230.285 76.590 230.550 77.600 ;
        RECT 234.125 77.025 234.475 78.275 ;
        RECT 236.240 77.850 237.450 78.370 ;
        RECT 237.620 77.680 238.830 78.200 ;
        RECT 239.920 77.850 241.130 78.370 ;
        RECT 230.720 76.590 236.065 77.025 ;
        RECT 236.240 76.590 238.830 77.680 ;
        RECT 239.460 76.590 239.750 77.755 ;
        RECT 241.300 77.680 242.510 78.200 ;
        RECT 243.615 78.150 243.835 78.550 ;
        RECT 242.680 77.950 243.170 78.150 ;
        RECT 243.360 77.940 243.835 78.150 ;
        RECT 244.080 78.150 244.290 78.550 ;
        RECT 244.545 78.485 245.300 78.610 ;
        RECT 244.545 78.440 245.390 78.485 ;
        RECT 245.120 78.320 245.390 78.440 ;
        RECT 244.080 77.940 244.410 78.150 ;
        RECT 244.580 77.880 244.990 78.185 ;
        RECT 239.920 76.590 242.510 77.680 ;
        RECT 242.685 77.710 243.860 77.770 ;
        RECT 245.220 77.745 245.390 78.320 ;
        RECT 245.190 77.710 245.390 77.745 ;
        RECT 242.685 77.600 245.390 77.710 ;
        RECT 242.685 76.980 242.940 77.600 ;
        RECT 243.530 77.540 245.330 77.600 ;
        RECT 243.530 77.510 243.860 77.540 ;
        RECT 245.560 77.440 245.730 78.640 ;
        RECT 246.440 78.570 246.610 78.920 ;
        RECT 246.810 78.740 247.140 79.140 ;
        RECT 247.310 78.570 247.480 78.920 ;
        RECT 247.650 78.740 248.030 79.140 ;
        RECT 245.905 77.900 246.255 78.470 ;
        RECT 246.440 78.400 248.050 78.570 ;
        RECT 248.220 78.465 248.490 78.810 ;
        RECT 248.660 78.595 254.005 79.140 ;
        RECT 247.880 78.230 248.050 78.400 ;
        RECT 246.425 77.780 247.135 78.230 ;
        RECT 247.305 77.900 247.710 78.230 ;
        RECT 247.880 77.900 248.150 78.230 ;
        RECT 243.190 77.340 243.375 77.430 ;
        RECT 243.965 77.340 244.800 77.350 ;
        RECT 243.190 77.140 244.800 77.340 ;
        RECT 243.190 77.100 243.420 77.140 ;
        RECT 242.685 76.760 243.020 76.980 ;
        RECT 244.025 76.590 244.380 76.970 ;
        RECT 244.550 76.760 244.800 77.140 ;
        RECT 245.050 76.590 245.300 77.370 ;
        RECT 245.470 76.760 245.730 77.440 ;
        RECT 245.905 77.440 246.225 77.730 ;
        RECT 246.420 77.610 247.135 77.780 ;
        RECT 247.880 77.730 248.050 77.900 ;
        RECT 248.320 77.730 248.490 78.465 ;
        RECT 250.245 77.765 250.585 78.595 ;
        RECT 254.180 78.370 257.690 79.140 ;
        RECT 258.325 78.375 258.780 79.140 ;
        RECT 259.055 78.760 260.355 78.970 ;
        RECT 260.610 78.780 260.940 79.140 ;
        RECT 260.185 78.610 260.355 78.760 ;
        RECT 261.110 78.640 261.370 78.970 ;
        RECT 261.140 78.630 261.370 78.640 ;
        RECT 247.325 77.560 248.050 77.730 ;
        RECT 247.325 77.440 247.495 77.560 ;
        RECT 245.905 77.270 247.495 77.440 ;
        RECT 245.905 76.810 247.560 77.100 ;
        RECT 247.730 76.590 248.010 77.390 ;
        RECT 248.220 76.760 248.490 77.730 ;
        RECT 252.065 77.025 252.415 78.275 ;
        RECT 254.180 77.850 255.830 78.370 ;
        RECT 256.000 77.680 257.690 78.200 ;
        RECT 259.255 78.150 259.475 78.550 ;
        RECT 258.320 77.950 258.810 78.150 ;
        RECT 259.000 77.940 259.475 78.150 ;
        RECT 259.720 78.150 259.930 78.550 ;
        RECT 260.185 78.485 260.940 78.610 ;
        RECT 260.185 78.440 261.030 78.485 ;
        RECT 260.760 78.320 261.030 78.440 ;
        RECT 259.720 77.940 260.050 78.150 ;
        RECT 260.220 77.880 260.630 78.185 ;
        RECT 248.660 76.590 254.005 77.025 ;
        RECT 254.180 76.590 257.690 77.680 ;
        RECT 258.325 77.710 259.500 77.770 ;
        RECT 260.860 77.745 261.030 78.320 ;
        RECT 260.830 77.710 261.030 77.745 ;
        RECT 258.325 77.600 261.030 77.710 ;
        RECT 258.325 76.980 258.580 77.600 ;
        RECT 259.170 77.540 260.970 77.600 ;
        RECT 259.170 77.510 259.500 77.540 ;
        RECT 261.200 77.440 261.370 78.630 ;
        RECT 261.545 78.375 262.000 79.140 ;
        RECT 262.275 78.760 263.575 78.970 ;
        RECT 263.830 78.780 264.160 79.140 ;
        RECT 263.405 78.610 263.575 78.760 ;
        RECT 264.330 78.640 264.590 78.970 ;
        RECT 264.360 78.630 264.590 78.640 ;
        RECT 262.475 78.150 262.695 78.550 ;
        RECT 261.540 77.950 262.030 78.150 ;
        RECT 262.220 77.940 262.695 78.150 ;
        RECT 262.940 78.150 263.150 78.550 ;
        RECT 263.405 78.485 264.160 78.610 ;
        RECT 263.405 78.440 264.250 78.485 ;
        RECT 263.980 78.320 264.250 78.440 ;
        RECT 262.940 77.940 263.270 78.150 ;
        RECT 263.440 77.880 263.850 78.185 ;
        RECT 258.830 77.340 259.015 77.430 ;
        RECT 259.605 77.340 260.440 77.350 ;
        RECT 258.830 77.140 260.440 77.340 ;
        RECT 258.830 77.100 259.060 77.140 ;
        RECT 258.325 76.760 258.660 76.980 ;
        RECT 259.665 76.590 260.020 76.970 ;
        RECT 260.190 76.760 260.440 77.140 ;
        RECT 260.690 76.590 260.940 77.370 ;
        RECT 261.110 76.760 261.370 77.440 ;
        RECT 261.545 77.710 262.720 77.770 ;
        RECT 264.080 77.745 264.250 78.320 ;
        RECT 264.050 77.710 264.250 77.745 ;
        RECT 261.545 77.600 264.250 77.710 ;
        RECT 261.545 76.980 261.800 77.600 ;
        RECT 262.390 77.540 264.190 77.600 ;
        RECT 262.390 77.510 262.720 77.540 ;
        RECT 264.420 77.440 264.590 78.630 ;
        RECT 265.220 78.415 265.510 79.140 ;
        RECT 265.680 78.680 266.240 78.970 ;
        RECT 266.410 78.680 266.660 79.140 ;
        RECT 262.050 77.340 262.235 77.430 ;
        RECT 262.825 77.340 263.660 77.350 ;
        RECT 262.050 77.140 263.660 77.340 ;
        RECT 262.050 77.100 262.280 77.140 ;
        RECT 261.545 76.760 261.880 76.980 ;
        RECT 262.885 76.590 263.240 76.970 ;
        RECT 263.410 76.760 263.660 77.140 ;
        RECT 263.910 76.590 264.160 77.370 ;
        RECT 264.330 76.760 264.590 77.440 ;
        RECT 265.220 76.590 265.510 77.755 ;
        RECT 265.680 77.310 265.930 78.680 ;
        RECT 267.280 78.510 267.610 78.870 ;
        RECT 267.980 78.595 273.325 79.140 ;
        RECT 273.500 78.595 278.845 79.140 ;
        RECT 266.220 78.320 267.610 78.510 ;
        RECT 266.220 78.230 266.390 78.320 ;
        RECT 266.100 77.900 266.390 78.230 ;
        RECT 266.560 77.900 266.900 78.150 ;
        RECT 267.120 77.900 267.795 78.150 ;
        RECT 266.220 77.650 266.390 77.900 ;
        RECT 266.220 77.480 267.160 77.650 ;
        RECT 267.530 77.540 267.795 77.900 ;
        RECT 269.565 77.765 269.905 78.595 ;
        RECT 265.680 76.760 266.140 77.310 ;
        RECT 266.330 76.590 266.660 77.310 ;
        RECT 266.860 76.930 267.160 77.480 ;
        RECT 267.330 76.590 267.610 77.260 ;
        RECT 271.385 77.025 271.735 78.275 ;
        RECT 275.085 77.765 275.425 78.595 ;
        RECT 279.945 78.430 280.200 78.960 ;
        RECT 280.370 78.680 280.675 79.140 ;
        RECT 280.920 78.760 281.990 78.930 ;
        RECT 276.905 77.025 277.255 78.275 ;
        RECT 279.945 77.780 280.155 78.430 ;
        RECT 280.920 78.405 281.240 78.760 ;
        RECT 280.915 78.230 281.240 78.405 ;
        RECT 280.325 77.930 281.240 78.230 ;
        RECT 281.410 78.190 281.650 78.590 ;
        RECT 281.820 78.530 281.990 78.760 ;
        RECT 282.160 78.700 282.350 79.140 ;
        RECT 282.520 78.690 283.470 78.970 ;
        RECT 283.690 78.780 284.040 78.950 ;
        RECT 281.820 78.360 282.350 78.530 ;
        RECT 280.325 77.900 281.065 77.930 ;
        RECT 267.980 76.590 273.325 77.025 ;
        RECT 273.500 76.590 278.845 77.025 ;
        RECT 279.945 76.900 280.200 77.780 ;
        RECT 280.370 76.590 280.675 77.730 ;
        RECT 280.895 77.310 281.065 77.900 ;
        RECT 281.410 77.820 281.950 78.190 ;
        RECT 282.130 78.080 282.350 78.360 ;
        RECT 282.520 77.910 282.690 78.690 ;
        RECT 282.285 77.740 282.690 77.910 ;
        RECT 282.860 77.900 283.210 78.520 ;
        RECT 282.285 77.650 282.455 77.740 ;
        RECT 283.380 77.730 283.590 78.520 ;
        RECT 281.235 77.480 282.455 77.650 ;
        RECT 282.915 77.570 283.590 77.730 ;
        RECT 280.895 77.140 281.695 77.310 ;
        RECT 281.015 76.590 281.345 76.970 ;
        RECT 281.525 76.850 281.695 77.140 ;
        RECT 282.285 77.100 282.455 77.480 ;
        RECT 282.625 77.560 283.590 77.570 ;
        RECT 283.780 78.390 284.040 78.780 ;
        RECT 284.250 78.680 284.580 79.140 ;
        RECT 285.455 78.750 286.310 78.920 ;
        RECT 286.515 78.750 287.010 78.920 ;
        RECT 287.180 78.780 287.510 79.140 ;
        RECT 283.780 77.700 283.950 78.390 ;
        RECT 284.120 78.040 284.290 78.220 ;
        RECT 284.460 78.210 285.250 78.460 ;
        RECT 285.455 78.040 285.625 78.750 ;
        RECT 285.795 78.240 286.150 78.460 ;
        RECT 284.120 77.870 285.810 78.040 ;
        RECT 282.625 77.270 283.085 77.560 ;
        RECT 283.780 77.530 285.280 77.700 ;
        RECT 283.780 77.390 283.950 77.530 ;
        RECT 283.390 77.220 283.950 77.390 ;
        RECT 281.865 76.590 282.115 77.050 ;
        RECT 282.285 76.760 283.155 77.100 ;
        RECT 283.390 76.760 283.560 77.220 ;
        RECT 284.395 77.190 285.470 77.360 ;
        RECT 283.730 76.590 284.100 77.050 ;
        RECT 284.395 76.850 284.565 77.190 ;
        RECT 284.735 76.590 285.065 77.020 ;
        RECT 285.300 76.850 285.470 77.190 ;
        RECT 285.640 77.090 285.810 77.870 ;
        RECT 285.980 77.650 286.150 78.240 ;
        RECT 286.320 77.840 286.670 78.460 ;
        RECT 285.980 77.260 286.445 77.650 ;
        RECT 286.840 77.390 287.010 78.750 ;
        RECT 287.180 77.560 287.640 78.610 ;
        RECT 286.615 77.220 287.010 77.390 ;
        RECT 286.615 77.090 286.785 77.220 ;
        RECT 285.640 76.760 286.320 77.090 ;
        RECT 286.535 76.760 286.785 77.090 ;
        RECT 286.955 76.590 287.205 77.050 ;
        RECT 287.375 76.775 287.700 77.560 ;
        RECT 287.870 76.760 288.040 78.880 ;
        RECT 288.210 78.760 288.540 79.140 ;
        RECT 288.710 78.590 288.965 78.880 ;
        RECT 288.215 78.420 288.965 78.590 ;
        RECT 288.215 77.430 288.445 78.420 ;
        RECT 289.140 78.370 290.810 79.140 ;
        RECT 290.980 78.415 291.270 79.140 ;
        RECT 291.500 78.680 291.745 79.140 ;
        RECT 288.615 77.600 288.965 78.250 ;
        RECT 289.140 77.850 289.890 78.370 ;
        RECT 290.060 77.680 290.810 78.200 ;
        RECT 291.440 77.900 291.755 78.510 ;
        RECT 291.925 78.150 292.175 78.960 ;
        RECT 292.345 78.615 292.605 79.140 ;
        RECT 292.775 78.490 293.035 78.945 ;
        RECT 293.205 78.660 293.465 79.140 ;
        RECT 293.635 78.490 293.895 78.945 ;
        RECT 294.065 78.660 294.325 79.140 ;
        RECT 294.495 78.490 294.755 78.945 ;
        RECT 294.925 78.660 295.185 79.140 ;
        RECT 295.355 78.490 295.615 78.945 ;
        RECT 295.785 78.660 296.085 79.140 ;
        RECT 292.775 78.320 296.085 78.490 ;
        RECT 291.925 77.900 294.945 78.150 ;
        RECT 288.215 77.260 288.965 77.430 ;
        RECT 288.210 76.590 288.540 77.090 ;
        RECT 288.710 76.760 288.965 77.260 ;
        RECT 289.140 76.590 290.810 77.680 ;
        RECT 290.980 76.590 291.270 77.755 ;
        RECT 291.450 76.590 291.745 77.700 ;
        RECT 291.925 76.765 292.175 77.900 ;
        RECT 295.115 77.730 296.085 78.320 ;
        RECT 296.500 78.390 297.710 79.140 ;
        RECT 297.885 78.590 298.140 78.880 ;
        RECT 298.310 78.760 298.640 79.140 ;
        RECT 297.885 78.420 298.635 78.590 ;
        RECT 296.500 77.850 297.020 78.390 ;
        RECT 292.345 76.590 292.605 77.700 ;
        RECT 292.775 77.490 296.085 77.730 ;
        RECT 297.190 77.680 297.710 78.220 ;
        RECT 292.775 76.765 293.035 77.490 ;
        RECT 293.205 76.590 293.465 77.320 ;
        RECT 293.635 76.765 293.895 77.490 ;
        RECT 294.065 76.590 294.325 77.320 ;
        RECT 294.495 76.765 294.755 77.490 ;
        RECT 294.925 76.590 295.185 77.320 ;
        RECT 295.355 76.765 295.615 77.490 ;
        RECT 295.785 76.590 296.080 77.320 ;
        RECT 296.500 76.590 297.710 77.680 ;
        RECT 297.885 77.600 298.235 78.250 ;
        RECT 298.405 77.430 298.635 78.420 ;
        RECT 297.885 77.260 298.635 77.430 ;
        RECT 297.885 76.760 298.140 77.260 ;
        RECT 298.310 76.590 298.640 77.090 ;
        RECT 298.810 76.760 298.980 78.880 ;
        RECT 299.340 78.780 299.670 79.140 ;
        RECT 299.840 78.750 300.335 78.920 ;
        RECT 300.540 78.750 301.395 78.920 ;
        RECT 299.210 77.560 299.670 78.610 ;
        RECT 299.150 76.775 299.475 77.560 ;
        RECT 299.840 77.390 300.010 78.750 ;
        RECT 300.180 77.840 300.530 78.460 ;
        RECT 300.700 78.240 301.055 78.460 ;
        RECT 300.700 77.650 300.870 78.240 ;
        RECT 301.225 78.040 301.395 78.750 ;
        RECT 302.270 78.680 302.600 79.140 ;
        RECT 302.810 78.780 303.160 78.950 ;
        RECT 301.600 78.210 302.390 78.460 ;
        RECT 302.810 78.390 303.070 78.780 ;
        RECT 303.380 78.690 304.330 78.970 ;
        RECT 304.500 78.700 304.690 79.140 ;
        RECT 304.860 78.760 305.930 78.930 ;
        RECT 302.560 78.040 302.730 78.220 ;
        RECT 299.840 77.220 300.235 77.390 ;
        RECT 300.405 77.260 300.870 77.650 ;
        RECT 301.040 77.870 302.730 78.040 ;
        RECT 300.065 77.090 300.235 77.220 ;
        RECT 301.040 77.090 301.210 77.870 ;
        RECT 302.900 77.700 303.070 78.390 ;
        RECT 301.570 77.530 303.070 77.700 ;
        RECT 303.260 77.730 303.470 78.520 ;
        RECT 303.640 77.900 303.990 78.520 ;
        RECT 304.160 77.910 304.330 78.690 ;
        RECT 304.860 78.530 305.030 78.760 ;
        RECT 304.500 78.360 305.030 78.530 ;
        RECT 304.500 78.080 304.720 78.360 ;
        RECT 305.200 78.190 305.440 78.590 ;
        RECT 304.160 77.740 304.565 77.910 ;
        RECT 304.900 77.820 305.440 78.190 ;
        RECT 305.610 78.405 305.930 78.760 ;
        RECT 306.175 78.680 306.480 79.140 ;
        RECT 306.650 78.430 306.900 78.960 ;
        RECT 305.610 78.230 305.935 78.405 ;
        RECT 305.610 77.930 306.525 78.230 ;
        RECT 305.785 77.900 306.525 77.930 ;
        RECT 303.260 77.570 303.935 77.730 ;
        RECT 304.395 77.650 304.565 77.740 ;
        RECT 303.260 77.560 304.225 77.570 ;
        RECT 302.900 77.390 303.070 77.530 ;
        RECT 299.645 76.590 299.895 77.050 ;
        RECT 300.065 76.760 300.315 77.090 ;
        RECT 300.530 76.760 301.210 77.090 ;
        RECT 301.380 77.190 302.455 77.360 ;
        RECT 302.900 77.220 303.460 77.390 ;
        RECT 303.765 77.270 304.225 77.560 ;
        RECT 304.395 77.480 305.615 77.650 ;
        RECT 301.380 76.850 301.550 77.190 ;
        RECT 301.785 76.590 302.115 77.020 ;
        RECT 302.285 76.850 302.455 77.190 ;
        RECT 302.750 76.590 303.120 77.050 ;
        RECT 303.290 76.760 303.460 77.220 ;
        RECT 304.395 77.100 304.565 77.480 ;
        RECT 305.785 77.310 305.955 77.900 ;
        RECT 306.695 77.780 306.900 78.430 ;
        RECT 307.070 78.385 307.320 79.140 ;
        RECT 307.540 78.370 309.210 79.140 ;
        RECT 309.840 78.390 311.050 79.140 ;
        RECT 307.540 77.850 308.290 78.370 ;
        RECT 303.695 76.760 304.565 77.100 ;
        RECT 305.155 77.140 305.955 77.310 ;
        RECT 304.735 76.590 304.985 77.050 ;
        RECT 305.155 76.850 305.325 77.140 ;
        RECT 305.505 76.590 305.835 76.970 ;
        RECT 306.175 76.590 306.480 77.730 ;
        RECT 306.650 76.900 306.900 77.780 ;
        RECT 307.070 76.590 307.320 77.730 ;
        RECT 308.460 77.680 309.210 78.200 ;
        RECT 307.540 76.590 309.210 77.680 ;
        RECT 309.840 77.680 310.360 78.220 ;
        RECT 310.530 77.850 311.050 78.390 ;
        RECT 309.840 76.590 311.050 77.680 ;
        RECT 162.095 76.420 311.135 76.590 ;
        RECT 162.180 75.330 163.390 76.420 ;
        RECT 163.560 75.330 165.230 76.420 ;
        RECT 165.865 75.750 166.120 76.250 ;
        RECT 166.290 75.920 166.620 76.420 ;
        RECT 165.865 75.580 166.615 75.750 ;
        RECT 162.180 74.620 162.700 75.160 ;
        RECT 162.870 74.790 163.390 75.330 ;
        RECT 163.560 74.640 164.310 75.160 ;
        RECT 164.480 74.810 165.230 75.330 ;
        RECT 165.865 74.760 166.215 75.410 ;
        RECT 162.180 73.870 163.390 74.620 ;
        RECT 163.560 73.870 165.230 74.640 ;
        RECT 166.385 74.590 166.615 75.580 ;
        RECT 165.865 74.420 166.615 74.590 ;
        RECT 165.865 74.130 166.120 74.420 ;
        RECT 166.290 73.870 166.620 74.250 ;
        RECT 166.790 74.130 166.960 76.250 ;
        RECT 167.130 75.450 167.455 76.235 ;
        RECT 167.625 75.960 167.875 76.420 ;
        RECT 168.045 75.920 168.295 76.250 ;
        RECT 168.510 75.920 169.190 76.250 ;
        RECT 168.045 75.790 168.215 75.920 ;
        RECT 167.820 75.620 168.215 75.790 ;
        RECT 167.190 74.400 167.650 75.450 ;
        RECT 167.820 74.260 167.990 75.620 ;
        RECT 168.385 75.360 168.850 75.750 ;
        RECT 168.160 74.550 168.510 75.170 ;
        RECT 168.680 74.770 168.850 75.360 ;
        RECT 169.020 75.140 169.190 75.920 ;
        RECT 169.360 75.820 169.530 76.160 ;
        RECT 169.765 75.990 170.095 76.420 ;
        RECT 170.265 75.820 170.435 76.160 ;
        RECT 170.730 75.960 171.100 76.420 ;
        RECT 169.360 75.650 170.435 75.820 ;
        RECT 171.270 75.790 171.440 76.250 ;
        RECT 171.675 75.910 172.545 76.250 ;
        RECT 172.715 75.960 172.965 76.420 ;
        RECT 170.880 75.620 171.440 75.790 ;
        RECT 170.880 75.480 171.050 75.620 ;
        RECT 169.550 75.310 171.050 75.480 ;
        RECT 171.745 75.450 172.205 75.740 ;
        RECT 169.020 74.970 170.710 75.140 ;
        RECT 168.680 74.550 169.035 74.770 ;
        RECT 169.205 74.260 169.375 74.970 ;
        RECT 169.580 74.550 170.370 74.800 ;
        RECT 170.540 74.790 170.710 74.970 ;
        RECT 170.880 74.620 171.050 75.310 ;
        RECT 167.320 73.870 167.650 74.230 ;
        RECT 167.820 74.090 168.315 74.260 ;
        RECT 168.520 74.090 169.375 74.260 ;
        RECT 170.250 73.870 170.580 74.330 ;
        RECT 170.790 74.230 171.050 74.620 ;
        RECT 171.240 75.440 172.205 75.450 ;
        RECT 172.375 75.530 172.545 75.910 ;
        RECT 173.135 75.870 173.305 76.160 ;
        RECT 173.485 76.040 173.815 76.420 ;
        RECT 173.135 75.700 173.935 75.870 ;
        RECT 171.240 75.280 171.915 75.440 ;
        RECT 172.375 75.360 173.595 75.530 ;
        RECT 171.240 74.490 171.450 75.280 ;
        RECT 172.375 75.270 172.545 75.360 ;
        RECT 171.620 74.490 171.970 75.110 ;
        RECT 172.140 75.100 172.545 75.270 ;
        RECT 172.140 74.320 172.310 75.100 ;
        RECT 172.480 74.650 172.700 74.930 ;
        RECT 172.880 74.820 173.420 75.190 ;
        RECT 173.765 75.110 173.935 75.700 ;
        RECT 174.155 75.280 174.460 76.420 ;
        RECT 174.630 75.230 174.885 76.110 ;
        RECT 175.060 75.255 175.350 76.420 ;
        RECT 175.525 75.280 175.860 76.250 ;
        RECT 176.030 75.280 176.200 76.420 ;
        RECT 176.370 76.080 178.400 76.250 ;
        RECT 173.765 75.080 174.505 75.110 ;
        RECT 172.480 74.480 173.010 74.650 ;
        RECT 170.790 74.060 171.140 74.230 ;
        RECT 171.360 74.040 172.310 74.320 ;
        RECT 172.480 73.870 172.670 74.310 ;
        RECT 172.840 74.250 173.010 74.480 ;
        RECT 173.180 74.420 173.420 74.820 ;
        RECT 173.590 74.780 174.505 75.080 ;
        RECT 173.590 74.605 173.915 74.780 ;
        RECT 173.590 74.250 173.910 74.605 ;
        RECT 174.675 74.580 174.885 75.230 ;
        RECT 175.525 74.610 175.695 75.280 ;
        RECT 176.370 75.110 176.540 76.080 ;
        RECT 175.865 74.780 176.120 75.110 ;
        RECT 176.345 74.780 176.540 75.110 ;
        RECT 176.710 75.740 177.835 75.910 ;
        RECT 175.950 74.610 176.120 74.780 ;
        RECT 176.710 74.610 176.880 75.740 ;
        RECT 172.840 74.080 173.910 74.250 ;
        RECT 174.155 73.870 174.460 74.330 ;
        RECT 174.630 74.050 174.885 74.580 ;
        RECT 175.060 73.870 175.350 74.595 ;
        RECT 175.525 74.040 175.780 74.610 ;
        RECT 175.950 74.440 176.880 74.610 ;
        RECT 177.050 75.400 178.060 75.570 ;
        RECT 177.050 74.600 177.220 75.400 ;
        RECT 176.705 74.405 176.880 74.440 ;
        RECT 175.950 73.870 176.280 74.270 ;
        RECT 176.705 74.040 177.235 74.405 ;
        RECT 177.425 74.380 177.700 75.200 ;
        RECT 177.420 74.210 177.700 74.380 ;
        RECT 177.425 74.040 177.700 74.210 ;
        RECT 177.870 74.040 178.060 75.400 ;
        RECT 178.230 75.415 178.400 76.080 ;
        RECT 178.570 75.660 178.740 76.420 ;
        RECT 178.975 75.660 179.490 76.070 ;
        RECT 178.230 75.225 178.980 75.415 ;
        RECT 179.150 74.850 179.490 75.660 ;
        RECT 179.660 75.330 180.870 76.420 ;
        RECT 181.045 75.750 181.300 76.250 ;
        RECT 181.470 75.920 181.800 76.420 ;
        RECT 181.045 75.580 181.795 75.750 ;
        RECT 178.260 74.680 179.490 74.850 ;
        RECT 178.240 73.870 178.750 74.405 ;
        RECT 178.970 74.075 179.215 74.680 ;
        RECT 179.660 74.620 180.180 75.160 ;
        RECT 180.350 74.790 180.870 75.330 ;
        RECT 181.045 74.760 181.395 75.410 ;
        RECT 179.660 73.870 180.870 74.620 ;
        RECT 181.565 74.590 181.795 75.580 ;
        RECT 181.045 74.420 181.795 74.590 ;
        RECT 181.045 74.130 181.300 74.420 ;
        RECT 181.470 73.870 181.800 74.250 ;
        RECT 181.970 74.130 182.140 76.250 ;
        RECT 182.310 75.450 182.635 76.235 ;
        RECT 182.805 75.960 183.055 76.420 ;
        RECT 183.225 75.920 183.475 76.250 ;
        RECT 183.690 75.920 184.370 76.250 ;
        RECT 183.225 75.790 183.395 75.920 ;
        RECT 183.000 75.620 183.395 75.790 ;
        RECT 182.370 74.400 182.830 75.450 ;
        RECT 183.000 74.260 183.170 75.620 ;
        RECT 183.565 75.360 184.030 75.750 ;
        RECT 183.340 74.550 183.690 75.170 ;
        RECT 183.860 74.770 184.030 75.360 ;
        RECT 184.200 75.140 184.370 75.920 ;
        RECT 184.540 75.820 184.710 76.160 ;
        RECT 184.945 75.990 185.275 76.420 ;
        RECT 185.445 75.820 185.615 76.160 ;
        RECT 185.910 75.960 186.280 76.420 ;
        RECT 184.540 75.650 185.615 75.820 ;
        RECT 186.450 75.790 186.620 76.250 ;
        RECT 186.855 75.910 187.725 76.250 ;
        RECT 187.895 75.960 188.145 76.420 ;
        RECT 186.060 75.620 186.620 75.790 ;
        RECT 186.060 75.480 186.230 75.620 ;
        RECT 184.730 75.310 186.230 75.480 ;
        RECT 186.925 75.450 187.385 75.740 ;
        RECT 184.200 74.970 185.890 75.140 ;
        RECT 183.860 74.550 184.215 74.770 ;
        RECT 184.385 74.260 184.555 74.970 ;
        RECT 184.760 74.550 185.550 74.800 ;
        RECT 185.720 74.790 185.890 74.970 ;
        RECT 186.060 74.620 186.230 75.310 ;
        RECT 182.500 73.870 182.830 74.230 ;
        RECT 183.000 74.090 183.495 74.260 ;
        RECT 183.700 74.090 184.555 74.260 ;
        RECT 185.430 73.870 185.760 74.330 ;
        RECT 185.970 74.230 186.230 74.620 ;
        RECT 186.420 75.440 187.385 75.450 ;
        RECT 187.555 75.530 187.725 75.910 ;
        RECT 188.315 75.870 188.485 76.160 ;
        RECT 188.665 76.040 188.995 76.420 ;
        RECT 188.315 75.700 189.115 75.870 ;
        RECT 186.420 75.280 187.095 75.440 ;
        RECT 187.555 75.360 188.775 75.530 ;
        RECT 186.420 74.490 186.630 75.280 ;
        RECT 187.555 75.270 187.725 75.360 ;
        RECT 186.800 74.490 187.150 75.110 ;
        RECT 187.320 75.100 187.725 75.270 ;
        RECT 187.320 74.320 187.490 75.100 ;
        RECT 187.660 74.650 187.880 74.930 ;
        RECT 188.060 74.820 188.600 75.190 ;
        RECT 188.945 75.110 189.115 75.700 ;
        RECT 189.335 75.280 189.640 76.420 ;
        RECT 189.810 75.230 190.065 76.110 ;
        RECT 190.240 75.330 191.450 76.420 ;
        RECT 191.625 75.750 191.880 76.250 ;
        RECT 192.050 75.920 192.380 76.420 ;
        RECT 191.625 75.580 192.375 75.750 ;
        RECT 188.945 75.080 189.685 75.110 ;
        RECT 187.660 74.480 188.190 74.650 ;
        RECT 185.970 74.060 186.320 74.230 ;
        RECT 186.540 74.040 187.490 74.320 ;
        RECT 187.660 73.870 187.850 74.310 ;
        RECT 188.020 74.250 188.190 74.480 ;
        RECT 188.360 74.420 188.600 74.820 ;
        RECT 188.770 74.780 189.685 75.080 ;
        RECT 188.770 74.605 189.095 74.780 ;
        RECT 188.770 74.250 189.090 74.605 ;
        RECT 189.855 74.580 190.065 75.230 ;
        RECT 188.020 74.080 189.090 74.250 ;
        RECT 189.335 73.870 189.640 74.330 ;
        RECT 189.810 74.050 190.065 74.580 ;
        RECT 190.240 74.620 190.760 75.160 ;
        RECT 190.930 74.790 191.450 75.330 ;
        RECT 191.625 74.760 191.975 75.410 ;
        RECT 190.240 73.870 191.450 74.620 ;
        RECT 192.145 74.590 192.375 75.580 ;
        RECT 191.625 74.420 192.375 74.590 ;
        RECT 191.625 74.130 191.880 74.420 ;
        RECT 192.050 73.870 192.380 74.250 ;
        RECT 192.550 74.130 192.720 76.250 ;
        RECT 192.890 75.450 193.215 76.235 ;
        RECT 193.385 75.960 193.635 76.420 ;
        RECT 193.805 75.920 194.055 76.250 ;
        RECT 194.270 75.920 194.950 76.250 ;
        RECT 193.805 75.790 193.975 75.920 ;
        RECT 193.580 75.620 193.975 75.790 ;
        RECT 192.950 74.400 193.410 75.450 ;
        RECT 193.580 74.260 193.750 75.620 ;
        RECT 194.145 75.360 194.610 75.750 ;
        RECT 193.920 74.550 194.270 75.170 ;
        RECT 194.440 74.770 194.610 75.360 ;
        RECT 194.780 75.140 194.950 75.920 ;
        RECT 195.120 75.820 195.290 76.160 ;
        RECT 195.525 75.990 195.855 76.420 ;
        RECT 196.025 75.820 196.195 76.160 ;
        RECT 196.490 75.960 196.860 76.420 ;
        RECT 195.120 75.650 196.195 75.820 ;
        RECT 197.030 75.790 197.200 76.250 ;
        RECT 197.435 75.910 198.305 76.250 ;
        RECT 198.475 75.960 198.725 76.420 ;
        RECT 196.640 75.620 197.200 75.790 ;
        RECT 196.640 75.480 196.810 75.620 ;
        RECT 195.310 75.310 196.810 75.480 ;
        RECT 197.505 75.450 197.965 75.740 ;
        RECT 194.780 74.970 196.470 75.140 ;
        RECT 194.440 74.550 194.795 74.770 ;
        RECT 194.965 74.260 195.135 74.970 ;
        RECT 195.340 74.550 196.130 74.800 ;
        RECT 196.300 74.790 196.470 74.970 ;
        RECT 196.640 74.620 196.810 75.310 ;
        RECT 193.080 73.870 193.410 74.230 ;
        RECT 193.580 74.090 194.075 74.260 ;
        RECT 194.280 74.090 195.135 74.260 ;
        RECT 196.010 73.870 196.340 74.330 ;
        RECT 196.550 74.230 196.810 74.620 ;
        RECT 197.000 75.440 197.965 75.450 ;
        RECT 198.135 75.530 198.305 75.910 ;
        RECT 198.895 75.870 199.065 76.160 ;
        RECT 199.245 76.040 199.575 76.420 ;
        RECT 198.895 75.700 199.695 75.870 ;
        RECT 197.000 75.280 197.675 75.440 ;
        RECT 198.135 75.360 199.355 75.530 ;
        RECT 197.000 74.490 197.210 75.280 ;
        RECT 198.135 75.270 198.305 75.360 ;
        RECT 197.380 74.490 197.730 75.110 ;
        RECT 197.900 75.100 198.305 75.270 ;
        RECT 197.900 74.320 198.070 75.100 ;
        RECT 198.240 74.650 198.460 74.930 ;
        RECT 198.640 74.820 199.180 75.190 ;
        RECT 199.525 75.110 199.695 75.700 ;
        RECT 199.915 75.280 200.220 76.420 ;
        RECT 200.390 75.230 200.645 76.110 ;
        RECT 200.820 75.255 201.110 76.420 ;
        RECT 201.285 75.270 201.545 76.420 ;
        RECT 201.720 75.345 201.975 76.250 ;
        RECT 202.145 75.660 202.475 76.420 ;
        RECT 202.690 75.490 202.860 76.250 ;
        RECT 199.525 75.080 200.265 75.110 ;
        RECT 198.240 74.480 198.770 74.650 ;
        RECT 196.550 74.060 196.900 74.230 ;
        RECT 197.120 74.040 198.070 74.320 ;
        RECT 198.240 73.870 198.430 74.310 ;
        RECT 198.600 74.250 198.770 74.480 ;
        RECT 198.940 74.420 199.180 74.820 ;
        RECT 199.350 74.780 200.265 75.080 ;
        RECT 199.350 74.605 199.675 74.780 ;
        RECT 199.350 74.250 199.670 74.605 ;
        RECT 200.435 74.580 200.645 75.230 ;
        RECT 198.600 74.080 199.670 74.250 ;
        RECT 199.915 73.870 200.220 74.330 ;
        RECT 200.390 74.050 200.645 74.580 ;
        RECT 200.820 73.870 201.110 74.595 ;
        RECT 201.285 73.870 201.545 74.710 ;
        RECT 201.720 74.615 201.890 75.345 ;
        RECT 202.145 75.320 202.860 75.490 ;
        RECT 203.120 75.330 206.630 76.420 ;
        RECT 202.145 75.110 202.315 75.320 ;
        RECT 202.060 74.780 202.315 75.110 ;
        RECT 201.720 74.040 201.975 74.615 ;
        RECT 202.145 74.590 202.315 74.780 ;
        RECT 202.595 74.770 202.950 75.140 ;
        RECT 203.120 74.640 204.770 75.160 ;
        RECT 204.940 74.810 206.630 75.330 ;
        RECT 207.265 75.230 207.520 76.110 ;
        RECT 207.690 75.280 207.995 76.420 ;
        RECT 208.335 76.040 208.665 76.420 ;
        RECT 208.845 75.870 209.015 76.160 ;
        RECT 209.185 75.960 209.435 76.420 ;
        RECT 208.215 75.700 209.015 75.870 ;
        RECT 209.605 75.910 210.475 76.250 ;
        RECT 202.145 74.420 202.860 74.590 ;
        RECT 202.145 73.870 202.475 74.250 ;
        RECT 202.690 74.040 202.860 74.420 ;
        RECT 203.120 73.870 206.630 74.640 ;
        RECT 207.265 74.580 207.475 75.230 ;
        RECT 208.215 75.110 208.385 75.700 ;
        RECT 209.605 75.530 209.775 75.910 ;
        RECT 210.710 75.790 210.880 76.250 ;
        RECT 211.050 75.960 211.420 76.420 ;
        RECT 211.715 75.820 211.885 76.160 ;
        RECT 212.055 75.990 212.385 76.420 ;
        RECT 212.620 75.820 212.790 76.160 ;
        RECT 208.555 75.360 209.775 75.530 ;
        RECT 209.945 75.450 210.405 75.740 ;
        RECT 210.710 75.620 211.270 75.790 ;
        RECT 211.715 75.650 212.790 75.820 ;
        RECT 212.960 75.920 213.640 76.250 ;
        RECT 213.855 75.920 214.105 76.250 ;
        RECT 214.275 75.960 214.525 76.420 ;
        RECT 211.100 75.480 211.270 75.620 ;
        RECT 209.945 75.440 210.910 75.450 ;
        RECT 209.605 75.270 209.775 75.360 ;
        RECT 210.235 75.280 210.910 75.440 ;
        RECT 207.645 75.080 208.385 75.110 ;
        RECT 207.645 74.780 208.560 75.080 ;
        RECT 208.235 74.605 208.560 74.780 ;
        RECT 207.265 74.050 207.520 74.580 ;
        RECT 207.690 73.870 207.995 74.330 ;
        RECT 208.240 74.250 208.560 74.605 ;
        RECT 208.730 74.820 209.270 75.190 ;
        RECT 209.605 75.100 210.010 75.270 ;
        RECT 208.730 74.420 208.970 74.820 ;
        RECT 209.450 74.650 209.670 74.930 ;
        RECT 209.140 74.480 209.670 74.650 ;
        RECT 209.140 74.250 209.310 74.480 ;
        RECT 209.840 74.320 210.010 75.100 ;
        RECT 210.180 74.490 210.530 75.110 ;
        RECT 210.700 74.490 210.910 75.280 ;
        RECT 211.100 75.310 212.600 75.480 ;
        RECT 211.100 74.620 211.270 75.310 ;
        RECT 212.960 75.140 213.130 75.920 ;
        RECT 213.935 75.790 214.105 75.920 ;
        RECT 211.440 74.970 213.130 75.140 ;
        RECT 213.300 75.360 213.765 75.750 ;
        RECT 213.935 75.620 214.330 75.790 ;
        RECT 211.440 74.790 211.610 74.970 ;
        RECT 208.240 74.080 209.310 74.250 ;
        RECT 209.480 73.870 209.670 74.310 ;
        RECT 209.840 74.040 210.790 74.320 ;
        RECT 211.100 74.230 211.360 74.620 ;
        RECT 211.780 74.550 212.570 74.800 ;
        RECT 211.010 74.060 211.360 74.230 ;
        RECT 211.570 73.870 211.900 74.330 ;
        RECT 212.775 74.260 212.945 74.970 ;
        RECT 213.300 74.770 213.470 75.360 ;
        RECT 213.115 74.550 213.470 74.770 ;
        RECT 213.640 74.550 213.990 75.170 ;
        RECT 214.160 74.260 214.330 75.620 ;
        RECT 214.695 75.450 215.020 76.235 ;
        RECT 214.500 74.400 214.960 75.450 ;
        RECT 212.775 74.090 213.630 74.260 ;
        RECT 213.835 74.090 214.330 74.260 ;
        RECT 214.500 73.870 214.830 74.230 ;
        RECT 215.190 74.130 215.360 76.250 ;
        RECT 215.530 75.920 215.860 76.420 ;
        RECT 216.030 75.750 216.285 76.250 ;
        RECT 215.535 75.580 216.285 75.750 ;
        RECT 215.535 74.590 215.765 75.580 ;
        RECT 215.935 74.760 216.285 75.410 ;
        RECT 216.465 75.280 216.800 76.250 ;
        RECT 216.970 75.280 217.140 76.420 ;
        RECT 217.310 76.080 219.340 76.250 ;
        RECT 216.465 74.610 216.635 75.280 ;
        RECT 217.310 75.110 217.480 76.080 ;
        RECT 216.805 74.780 217.060 75.110 ;
        RECT 217.285 74.780 217.480 75.110 ;
        RECT 217.650 75.740 218.775 75.910 ;
        RECT 216.890 74.610 217.060 74.780 ;
        RECT 217.650 74.610 217.820 75.740 ;
        RECT 215.535 74.420 216.285 74.590 ;
        RECT 215.530 73.870 215.860 74.250 ;
        RECT 216.030 74.130 216.285 74.420 ;
        RECT 216.465 74.040 216.720 74.610 ;
        RECT 216.890 74.440 217.820 74.610 ;
        RECT 217.990 75.400 219.000 75.570 ;
        RECT 217.990 74.600 218.160 75.400 ;
        RECT 217.645 74.405 217.820 74.440 ;
        RECT 216.890 73.870 217.220 74.270 ;
        RECT 217.645 74.040 218.175 74.405 ;
        RECT 218.365 74.380 218.640 75.200 ;
        RECT 218.360 74.210 218.640 74.380 ;
        RECT 218.365 74.040 218.640 74.210 ;
        RECT 218.810 74.040 219.000 75.400 ;
        RECT 219.170 75.415 219.340 76.080 ;
        RECT 219.510 75.660 219.680 76.420 ;
        RECT 219.915 75.660 220.430 76.070 ;
        RECT 219.170 75.225 219.920 75.415 ;
        RECT 220.090 74.850 220.430 75.660 ;
        RECT 220.600 75.330 223.190 76.420 ;
        RECT 219.200 74.680 220.430 74.850 ;
        RECT 219.180 73.870 219.690 74.405 ;
        RECT 219.910 74.075 220.155 74.680 ;
        RECT 220.600 74.640 221.810 75.160 ;
        RECT 221.980 74.810 223.190 75.330 ;
        RECT 223.825 75.270 224.085 76.420 ;
        RECT 224.260 75.345 224.515 76.250 ;
        RECT 224.685 75.660 225.015 76.420 ;
        RECT 225.230 75.490 225.400 76.250 ;
        RECT 220.600 73.870 223.190 74.640 ;
        RECT 223.825 73.870 224.085 74.710 ;
        RECT 224.260 74.615 224.430 75.345 ;
        RECT 224.685 75.320 225.400 75.490 ;
        RECT 224.685 75.110 224.855 75.320 ;
        RECT 226.580 75.255 226.870 76.420 ;
        RECT 227.040 75.985 232.385 76.420 ;
        RECT 232.560 75.985 237.905 76.420 ;
        RECT 238.080 75.985 243.425 76.420 ;
        RECT 243.600 75.985 248.945 76.420 ;
        RECT 224.600 74.780 224.855 75.110 ;
        RECT 224.260 74.040 224.515 74.615 ;
        RECT 224.685 74.590 224.855 74.780 ;
        RECT 225.135 74.770 225.490 75.140 ;
        RECT 224.685 74.420 225.400 74.590 ;
        RECT 224.685 73.870 225.015 74.250 ;
        RECT 225.230 74.040 225.400 74.420 ;
        RECT 226.580 73.870 226.870 74.595 ;
        RECT 228.625 74.415 228.965 75.245 ;
        RECT 230.445 74.735 230.795 75.985 ;
        RECT 234.145 74.415 234.485 75.245 ;
        RECT 235.965 74.735 236.315 75.985 ;
        RECT 239.665 74.415 240.005 75.245 ;
        RECT 241.485 74.735 241.835 75.985 ;
        RECT 245.185 74.415 245.525 75.245 ;
        RECT 247.005 74.735 247.355 75.985 ;
        RECT 249.120 75.330 251.710 76.420 ;
        RECT 249.120 74.640 250.330 75.160 ;
        RECT 250.500 74.810 251.710 75.330 ;
        RECT 252.340 75.255 252.630 76.420 ;
        RECT 252.800 75.985 258.145 76.420 ;
        RECT 227.040 73.870 232.385 74.415 ;
        RECT 232.560 73.870 237.905 74.415 ;
        RECT 238.080 73.870 243.425 74.415 ;
        RECT 243.600 73.870 248.945 74.415 ;
        RECT 249.120 73.870 251.710 74.640 ;
        RECT 252.340 73.870 252.630 74.595 ;
        RECT 254.385 74.415 254.725 75.245 ;
        RECT 256.205 74.735 256.555 75.985 ;
        RECT 258.320 75.330 259.990 76.420 ;
        RECT 258.320 74.640 259.070 75.160 ;
        RECT 259.240 74.810 259.990 75.330 ;
        RECT 260.250 75.410 260.420 76.250 ;
        RECT 260.590 76.080 261.760 76.250 ;
        RECT 260.590 75.580 260.920 76.080 ;
        RECT 261.430 76.040 261.760 76.080 ;
        RECT 261.950 76.000 262.305 76.420 ;
        RECT 261.090 75.820 261.320 75.910 ;
        RECT 262.475 75.820 262.725 76.250 ;
        RECT 261.090 75.580 262.725 75.820 ;
        RECT 262.895 75.660 263.225 76.420 ;
        RECT 263.395 75.580 263.650 76.250 ;
        RECT 263.840 75.985 269.185 76.420 ;
        RECT 269.360 75.985 274.705 76.420 ;
        RECT 260.250 75.240 263.310 75.410 ;
        RECT 260.165 74.860 260.515 75.070 ;
        RECT 260.685 74.860 261.130 75.060 ;
        RECT 261.300 74.860 261.775 75.060 ;
        RECT 252.800 73.870 258.145 74.415 ;
        RECT 258.320 73.870 259.990 74.640 ;
        RECT 260.250 74.520 261.315 74.690 ;
        RECT 260.250 74.040 260.420 74.520 ;
        RECT 260.590 73.870 260.920 74.350 ;
        RECT 261.145 74.290 261.315 74.520 ;
        RECT 261.495 74.460 261.775 74.860 ;
        RECT 262.045 74.860 262.375 75.060 ;
        RECT 262.545 74.890 262.920 75.060 ;
        RECT 262.545 74.860 262.910 74.890 ;
        RECT 262.045 74.460 262.330 74.860 ;
        RECT 263.140 74.690 263.310 75.240 ;
        RECT 262.510 74.520 263.310 74.690 ;
        RECT 262.510 74.290 262.680 74.520 ;
        RECT 263.480 74.450 263.650 75.580 ;
        RECT 263.465 74.380 263.650 74.450 ;
        RECT 265.425 74.415 265.765 75.245 ;
        RECT 267.245 74.735 267.595 75.985 ;
        RECT 270.945 74.415 271.285 75.245 ;
        RECT 272.765 74.735 273.115 75.985 ;
        RECT 274.900 75.570 275.230 76.420 ;
        RECT 275.400 76.080 276.510 76.250 ;
        RECT 275.400 75.570 275.620 76.080 ;
        RECT 276.320 75.920 276.510 76.080 ;
        RECT 276.705 75.960 277.035 76.420 ;
        RECT 275.790 75.750 276.090 75.910 ;
        RECT 277.205 75.750 277.440 76.250 ;
        RECT 275.790 75.570 277.440 75.750 ;
        RECT 274.915 75.230 276.890 75.400 ;
        RECT 274.915 74.840 275.245 75.230 ;
        RECT 275.415 74.860 276.215 75.060 ;
        RECT 276.395 74.860 276.890 75.230 ;
        RECT 274.900 74.500 277.060 74.670 ;
        RECT 263.440 74.370 263.650 74.380 ;
        RECT 261.145 74.040 262.680 74.290 ;
        RECT 262.850 73.870 263.180 74.350 ;
        RECT 263.395 74.040 263.650 74.370 ;
        RECT 263.840 73.870 269.185 74.415 ;
        RECT 269.360 73.870 274.705 74.415 ;
        RECT 274.900 74.040 275.230 74.500 ;
        RECT 275.410 73.870 275.580 74.330 ;
        RECT 275.760 74.040 276.090 74.500 ;
        RECT 276.320 73.870 276.490 74.330 ;
        RECT 276.730 74.210 277.060 74.500 ;
        RECT 277.230 74.380 277.440 75.570 ;
        RECT 277.610 75.355 277.920 76.420 ;
        RECT 278.100 75.255 278.390 76.420 ;
        RECT 279.025 75.230 279.280 76.110 ;
        RECT 279.450 75.280 279.755 76.420 ;
        RECT 280.095 76.040 280.425 76.420 ;
        RECT 280.605 75.870 280.775 76.160 ;
        RECT 280.945 75.960 281.195 76.420 ;
        RECT 279.975 75.700 280.775 75.870 ;
        RECT 281.365 75.910 282.235 76.250 ;
        RECT 277.610 74.550 277.925 75.185 ;
        RECT 277.610 74.210 277.920 74.380 ;
        RECT 276.730 74.040 277.920 74.210 ;
        RECT 278.100 73.870 278.390 74.595 ;
        RECT 279.025 74.580 279.235 75.230 ;
        RECT 279.975 75.110 280.145 75.700 ;
        RECT 281.365 75.530 281.535 75.910 ;
        RECT 282.470 75.790 282.640 76.250 ;
        RECT 282.810 75.960 283.180 76.420 ;
        RECT 283.475 75.820 283.645 76.160 ;
        RECT 283.815 75.990 284.145 76.420 ;
        RECT 284.380 75.820 284.550 76.160 ;
        RECT 280.315 75.360 281.535 75.530 ;
        RECT 281.705 75.450 282.165 75.740 ;
        RECT 282.470 75.620 283.030 75.790 ;
        RECT 283.475 75.650 284.550 75.820 ;
        RECT 284.720 75.920 285.400 76.250 ;
        RECT 285.615 75.920 285.865 76.250 ;
        RECT 286.035 75.960 286.285 76.420 ;
        RECT 282.860 75.480 283.030 75.620 ;
        RECT 281.705 75.440 282.670 75.450 ;
        RECT 281.365 75.270 281.535 75.360 ;
        RECT 281.995 75.280 282.670 75.440 ;
        RECT 279.405 75.080 280.145 75.110 ;
        RECT 279.405 74.780 280.320 75.080 ;
        RECT 279.995 74.605 280.320 74.780 ;
        RECT 279.025 74.050 279.280 74.580 ;
        RECT 279.450 73.870 279.755 74.330 ;
        RECT 280.000 74.250 280.320 74.605 ;
        RECT 280.490 74.820 281.030 75.190 ;
        RECT 281.365 75.100 281.770 75.270 ;
        RECT 280.490 74.420 280.730 74.820 ;
        RECT 281.210 74.650 281.430 74.930 ;
        RECT 280.900 74.480 281.430 74.650 ;
        RECT 280.900 74.250 281.070 74.480 ;
        RECT 281.600 74.320 281.770 75.100 ;
        RECT 281.940 74.490 282.290 75.110 ;
        RECT 282.460 74.490 282.670 75.280 ;
        RECT 282.860 75.310 284.360 75.480 ;
        RECT 282.860 74.620 283.030 75.310 ;
        RECT 284.720 75.140 284.890 75.920 ;
        RECT 285.695 75.790 285.865 75.920 ;
        RECT 283.200 74.970 284.890 75.140 ;
        RECT 285.060 75.360 285.525 75.750 ;
        RECT 285.695 75.620 286.090 75.790 ;
        RECT 283.200 74.790 283.370 74.970 ;
        RECT 280.000 74.080 281.070 74.250 ;
        RECT 281.240 73.870 281.430 74.310 ;
        RECT 281.600 74.040 282.550 74.320 ;
        RECT 282.860 74.230 283.120 74.620 ;
        RECT 283.540 74.550 284.330 74.800 ;
        RECT 282.770 74.060 283.120 74.230 ;
        RECT 283.330 73.870 283.660 74.330 ;
        RECT 284.535 74.260 284.705 74.970 ;
        RECT 285.060 74.770 285.230 75.360 ;
        RECT 284.875 74.550 285.230 74.770 ;
        RECT 285.400 74.550 285.750 75.170 ;
        RECT 285.920 74.260 286.090 75.620 ;
        RECT 286.455 75.450 286.780 76.235 ;
        RECT 286.260 74.400 286.720 75.450 ;
        RECT 284.535 74.090 285.390 74.260 ;
        RECT 285.595 74.090 286.090 74.260 ;
        RECT 286.260 73.870 286.590 74.230 ;
        RECT 286.950 74.130 287.120 76.250 ;
        RECT 287.290 75.920 287.620 76.420 ;
        RECT 287.790 75.750 288.045 76.250 ;
        RECT 287.295 75.580 288.045 75.750 ;
        RECT 287.295 74.590 287.525 75.580 ;
        RECT 287.695 74.760 288.045 75.410 ;
        RECT 288.220 75.330 289.430 76.420 ;
        RECT 288.220 74.620 288.740 75.160 ;
        RECT 288.910 74.790 289.430 75.330 ;
        RECT 289.610 75.310 289.905 76.420 ;
        RECT 290.085 75.110 290.335 76.245 ;
        RECT 290.505 75.310 290.765 76.420 ;
        RECT 290.935 75.520 291.195 76.245 ;
        RECT 291.365 75.690 291.625 76.420 ;
        RECT 291.795 75.520 292.055 76.245 ;
        RECT 292.225 75.690 292.485 76.420 ;
        RECT 292.655 75.520 292.915 76.245 ;
        RECT 293.085 75.690 293.345 76.420 ;
        RECT 293.515 75.520 293.775 76.245 ;
        RECT 293.945 75.690 294.240 76.420 ;
        RECT 294.665 75.750 294.920 76.250 ;
        RECT 295.090 75.920 295.420 76.420 ;
        RECT 294.665 75.580 295.415 75.750 ;
        RECT 290.935 75.280 294.245 75.520 ;
        RECT 287.295 74.420 288.045 74.590 ;
        RECT 287.290 73.870 287.620 74.250 ;
        RECT 287.790 74.130 288.045 74.420 ;
        RECT 288.220 73.870 289.430 74.620 ;
        RECT 289.600 74.500 289.915 75.110 ;
        RECT 290.085 74.860 293.105 75.110 ;
        RECT 289.660 73.870 289.905 74.330 ;
        RECT 290.085 74.050 290.335 74.860 ;
        RECT 293.275 74.690 294.245 75.280 ;
        RECT 294.665 74.760 295.015 75.410 ;
        RECT 290.935 74.520 294.245 74.690 ;
        RECT 295.185 74.590 295.415 75.580 ;
        RECT 290.505 73.870 290.765 74.395 ;
        RECT 290.935 74.065 291.195 74.520 ;
        RECT 291.365 73.870 291.625 74.350 ;
        RECT 291.795 74.065 292.055 74.520 ;
        RECT 292.225 73.870 292.485 74.350 ;
        RECT 292.655 74.065 292.915 74.520 ;
        RECT 293.085 73.870 293.345 74.350 ;
        RECT 293.515 74.065 293.775 74.520 ;
        RECT 294.665 74.420 295.415 74.590 ;
        RECT 293.945 73.870 294.245 74.350 ;
        RECT 294.665 74.130 294.920 74.420 ;
        RECT 295.090 73.870 295.420 74.250 ;
        RECT 295.590 74.130 295.760 76.250 ;
        RECT 295.930 75.450 296.255 76.235 ;
        RECT 296.425 75.960 296.675 76.420 ;
        RECT 296.845 75.920 297.095 76.250 ;
        RECT 297.310 75.920 297.990 76.250 ;
        RECT 296.845 75.790 297.015 75.920 ;
        RECT 296.620 75.620 297.015 75.790 ;
        RECT 295.990 74.400 296.450 75.450 ;
        RECT 296.620 74.260 296.790 75.620 ;
        RECT 297.185 75.360 297.650 75.750 ;
        RECT 296.960 74.550 297.310 75.170 ;
        RECT 297.480 74.770 297.650 75.360 ;
        RECT 297.820 75.140 297.990 75.920 ;
        RECT 298.160 75.820 298.330 76.160 ;
        RECT 298.565 75.990 298.895 76.420 ;
        RECT 299.065 75.820 299.235 76.160 ;
        RECT 299.530 75.960 299.900 76.420 ;
        RECT 298.160 75.650 299.235 75.820 ;
        RECT 300.070 75.790 300.240 76.250 ;
        RECT 300.475 75.910 301.345 76.250 ;
        RECT 301.515 75.960 301.765 76.420 ;
        RECT 299.680 75.620 300.240 75.790 ;
        RECT 299.680 75.480 299.850 75.620 ;
        RECT 298.350 75.310 299.850 75.480 ;
        RECT 300.545 75.450 301.005 75.740 ;
        RECT 297.820 74.970 299.510 75.140 ;
        RECT 297.480 74.550 297.835 74.770 ;
        RECT 298.005 74.260 298.175 74.970 ;
        RECT 298.380 74.550 299.170 74.800 ;
        RECT 299.340 74.790 299.510 74.970 ;
        RECT 299.680 74.620 299.850 75.310 ;
        RECT 296.120 73.870 296.450 74.230 ;
        RECT 296.620 74.090 297.115 74.260 ;
        RECT 297.320 74.090 298.175 74.260 ;
        RECT 299.050 73.870 299.380 74.330 ;
        RECT 299.590 74.230 299.850 74.620 ;
        RECT 300.040 75.440 301.005 75.450 ;
        RECT 301.175 75.530 301.345 75.910 ;
        RECT 301.935 75.870 302.105 76.160 ;
        RECT 302.285 76.040 302.615 76.420 ;
        RECT 301.935 75.700 302.735 75.870 ;
        RECT 300.040 75.280 300.715 75.440 ;
        RECT 301.175 75.360 302.395 75.530 ;
        RECT 300.040 74.490 300.250 75.280 ;
        RECT 301.175 75.270 301.345 75.360 ;
        RECT 300.420 74.490 300.770 75.110 ;
        RECT 300.940 75.100 301.345 75.270 ;
        RECT 300.940 74.320 301.110 75.100 ;
        RECT 301.280 74.650 301.500 74.930 ;
        RECT 301.680 74.820 302.220 75.190 ;
        RECT 302.565 75.110 302.735 75.700 ;
        RECT 302.955 75.280 303.260 76.420 ;
        RECT 303.430 75.230 303.685 76.110 ;
        RECT 303.860 75.255 304.150 76.420 ;
        RECT 304.325 75.280 304.660 76.250 ;
        RECT 304.830 75.280 305.000 76.420 ;
        RECT 305.170 76.080 307.200 76.250 ;
        RECT 302.565 75.080 303.305 75.110 ;
        RECT 301.280 74.480 301.810 74.650 ;
        RECT 299.590 74.060 299.940 74.230 ;
        RECT 300.160 74.040 301.110 74.320 ;
        RECT 301.280 73.870 301.470 74.310 ;
        RECT 301.640 74.250 301.810 74.480 ;
        RECT 301.980 74.420 302.220 74.820 ;
        RECT 302.390 74.780 303.305 75.080 ;
        RECT 302.390 74.605 302.715 74.780 ;
        RECT 302.390 74.250 302.710 74.605 ;
        RECT 303.475 74.580 303.685 75.230 ;
        RECT 304.325 74.610 304.495 75.280 ;
        RECT 305.170 75.110 305.340 76.080 ;
        RECT 304.665 74.780 304.920 75.110 ;
        RECT 305.145 74.780 305.340 75.110 ;
        RECT 305.510 75.740 306.635 75.910 ;
        RECT 304.750 74.610 304.920 74.780 ;
        RECT 305.510 74.610 305.680 75.740 ;
        RECT 301.640 74.080 302.710 74.250 ;
        RECT 302.955 73.870 303.260 74.330 ;
        RECT 303.430 74.050 303.685 74.580 ;
        RECT 303.860 73.870 304.150 74.595 ;
        RECT 304.325 74.040 304.580 74.610 ;
        RECT 304.750 74.440 305.680 74.610 ;
        RECT 305.850 75.400 306.860 75.570 ;
        RECT 305.850 74.600 306.020 75.400 ;
        RECT 306.225 75.060 306.500 75.200 ;
        RECT 306.220 74.890 306.500 75.060 ;
        RECT 305.505 74.405 305.680 74.440 ;
        RECT 304.750 73.870 305.080 74.270 ;
        RECT 305.505 74.040 306.035 74.405 ;
        RECT 306.225 74.040 306.500 74.890 ;
        RECT 306.670 74.040 306.860 75.400 ;
        RECT 307.030 75.415 307.200 76.080 ;
        RECT 307.370 75.660 307.540 76.420 ;
        RECT 307.775 75.660 308.290 76.070 ;
        RECT 307.030 75.225 307.780 75.415 ;
        RECT 307.950 74.850 308.290 75.660 ;
        RECT 308.460 75.330 309.670 76.420 ;
        RECT 307.060 74.680 308.290 74.850 ;
        RECT 307.040 73.870 307.550 74.405 ;
        RECT 307.770 74.075 308.015 74.680 ;
        RECT 308.460 74.620 308.980 75.160 ;
        RECT 309.150 74.790 309.670 75.330 ;
        RECT 309.840 75.330 311.050 76.420 ;
        RECT 309.840 74.790 310.360 75.330 ;
        RECT 310.530 74.620 311.050 75.160 ;
        RECT 308.460 73.870 309.670 74.620 ;
        RECT 309.840 73.870 311.050 74.620 ;
        RECT 162.095 73.700 311.135 73.870 ;
        RECT 162.180 72.950 163.390 73.700 ;
        RECT 163.560 73.155 168.905 73.700 ;
        RECT 162.180 72.410 162.700 72.950 ;
        RECT 162.870 72.240 163.390 72.780 ;
        RECT 165.145 72.325 165.485 73.155 ;
        RECT 170.005 73.150 170.260 73.440 ;
        RECT 170.430 73.320 170.760 73.700 ;
        RECT 170.005 72.980 170.755 73.150 ;
        RECT 162.180 71.150 163.390 72.240 ;
        RECT 166.965 71.585 167.315 72.835 ;
        RECT 170.005 72.160 170.355 72.810 ;
        RECT 170.525 71.990 170.755 72.980 ;
        RECT 170.005 71.820 170.755 71.990 ;
        RECT 163.560 71.150 168.905 71.585 ;
        RECT 170.005 71.320 170.260 71.820 ;
        RECT 170.430 71.150 170.760 71.650 ;
        RECT 170.930 71.320 171.100 73.440 ;
        RECT 171.460 73.340 171.790 73.700 ;
        RECT 171.960 73.310 172.455 73.480 ;
        RECT 172.660 73.310 173.515 73.480 ;
        RECT 171.330 72.120 171.790 73.170 ;
        RECT 171.270 71.335 171.595 72.120 ;
        RECT 171.960 71.950 172.130 73.310 ;
        RECT 172.300 72.400 172.650 73.020 ;
        RECT 172.820 72.800 173.175 73.020 ;
        RECT 172.820 72.210 172.990 72.800 ;
        RECT 173.345 72.600 173.515 73.310 ;
        RECT 174.390 73.240 174.720 73.700 ;
        RECT 174.930 73.340 175.280 73.510 ;
        RECT 173.720 72.770 174.510 73.020 ;
        RECT 174.930 72.950 175.190 73.340 ;
        RECT 175.500 73.250 176.450 73.530 ;
        RECT 176.620 73.260 176.810 73.700 ;
        RECT 176.980 73.320 178.050 73.490 ;
        RECT 174.680 72.600 174.850 72.780 ;
        RECT 171.960 71.780 172.355 71.950 ;
        RECT 172.525 71.820 172.990 72.210 ;
        RECT 173.160 72.430 174.850 72.600 ;
        RECT 172.185 71.650 172.355 71.780 ;
        RECT 173.160 71.650 173.330 72.430 ;
        RECT 175.020 72.260 175.190 72.950 ;
        RECT 173.690 72.090 175.190 72.260 ;
        RECT 175.380 72.290 175.590 73.080 ;
        RECT 175.760 72.460 176.110 73.080 ;
        RECT 176.280 72.470 176.450 73.250 ;
        RECT 176.980 73.090 177.150 73.320 ;
        RECT 176.620 72.920 177.150 73.090 ;
        RECT 176.620 72.640 176.840 72.920 ;
        RECT 177.320 72.750 177.560 73.150 ;
        RECT 176.280 72.300 176.685 72.470 ;
        RECT 177.020 72.380 177.560 72.750 ;
        RECT 177.730 72.965 178.050 73.320 ;
        RECT 178.295 73.240 178.600 73.700 ;
        RECT 178.770 72.990 179.020 73.520 ;
        RECT 177.730 72.790 178.055 72.965 ;
        RECT 177.730 72.490 178.645 72.790 ;
        RECT 177.905 72.460 178.645 72.490 ;
        RECT 175.380 72.130 176.055 72.290 ;
        RECT 176.515 72.210 176.685 72.300 ;
        RECT 175.380 72.120 176.345 72.130 ;
        RECT 175.020 71.950 175.190 72.090 ;
        RECT 171.765 71.150 172.015 71.610 ;
        RECT 172.185 71.320 172.435 71.650 ;
        RECT 172.650 71.320 173.330 71.650 ;
        RECT 173.500 71.750 174.575 71.920 ;
        RECT 175.020 71.780 175.580 71.950 ;
        RECT 175.885 71.830 176.345 72.120 ;
        RECT 176.515 72.040 177.735 72.210 ;
        RECT 173.500 71.410 173.670 71.750 ;
        RECT 173.905 71.150 174.235 71.580 ;
        RECT 174.405 71.410 174.575 71.750 ;
        RECT 174.870 71.150 175.240 71.610 ;
        RECT 175.410 71.320 175.580 71.780 ;
        RECT 176.515 71.660 176.685 72.040 ;
        RECT 177.905 71.870 178.075 72.460 ;
        RECT 178.815 72.340 179.020 72.990 ;
        RECT 179.190 72.945 179.440 73.700 ;
        RECT 179.660 72.930 183.170 73.700 ;
        RECT 183.340 72.950 184.550 73.700 ;
        RECT 184.820 73.235 185.070 73.700 ;
        RECT 185.240 73.060 185.410 73.530 ;
        RECT 185.660 73.240 185.830 73.700 ;
        RECT 186.080 73.060 186.250 73.530 ;
        RECT 186.500 73.240 186.670 73.700 ;
        RECT 186.920 73.060 187.090 73.530 ;
        RECT 187.460 73.240 187.725 73.700 ;
        RECT 179.660 72.410 181.310 72.930 ;
        RECT 175.815 71.320 176.685 71.660 ;
        RECT 177.275 71.700 178.075 71.870 ;
        RECT 176.855 71.150 177.105 71.610 ;
        RECT 177.275 71.410 177.445 71.700 ;
        RECT 177.625 71.150 177.955 71.530 ;
        RECT 178.295 71.150 178.600 72.290 ;
        RECT 178.770 71.460 179.020 72.340 ;
        RECT 179.190 71.150 179.440 72.290 ;
        RECT 181.480 72.240 183.170 72.760 ;
        RECT 183.340 72.410 183.860 72.950 ;
        RECT 184.720 72.880 187.090 73.060 ;
        RECT 187.940 72.975 188.230 73.700 ;
        RECT 189.105 73.220 189.405 73.700 ;
        RECT 189.575 73.050 189.835 73.505 ;
        RECT 190.005 73.220 190.265 73.700 ;
        RECT 190.435 73.050 190.695 73.505 ;
        RECT 190.865 73.220 191.125 73.700 ;
        RECT 191.295 73.050 191.555 73.505 ;
        RECT 191.725 73.220 191.985 73.700 ;
        RECT 192.155 73.050 192.415 73.505 ;
        RECT 192.585 73.175 192.845 73.700 ;
        RECT 189.105 72.880 192.415 73.050 ;
        RECT 184.030 72.240 184.550 72.780 ;
        RECT 179.660 71.150 183.170 72.240 ;
        RECT 183.340 71.150 184.550 72.240 ;
        RECT 184.720 72.290 185.070 72.880 ;
        RECT 185.240 72.460 187.750 72.710 ;
        RECT 184.720 72.120 187.170 72.290 ;
        RECT 184.720 72.100 185.490 72.120 ;
        RECT 184.820 71.150 184.990 71.610 ;
        RECT 185.160 71.320 185.490 72.100 ;
        RECT 185.660 71.150 185.830 71.950 ;
        RECT 186.000 71.320 186.330 72.120 ;
        RECT 186.500 71.150 186.670 71.950 ;
        RECT 186.840 71.320 187.170 72.120 ;
        RECT 187.430 71.150 187.725 72.290 ;
        RECT 187.940 71.150 188.230 72.315 ;
        RECT 189.105 72.290 190.075 72.880 ;
        RECT 193.015 72.710 193.265 73.520 ;
        RECT 193.445 73.240 193.690 73.700 ;
        RECT 190.245 72.460 193.265 72.710 ;
        RECT 193.435 72.460 193.750 73.070 ;
        RECT 193.920 72.930 196.510 73.700 ;
        RECT 196.685 72.960 196.940 73.530 ;
        RECT 197.110 73.300 197.440 73.700 ;
        RECT 197.865 73.165 198.395 73.530 ;
        RECT 197.865 73.130 198.040 73.165 ;
        RECT 197.110 72.960 198.040 73.130 ;
        RECT 198.585 73.020 198.860 73.530 ;
        RECT 189.105 72.050 192.415 72.290 ;
        RECT 189.110 71.150 189.405 71.880 ;
        RECT 189.575 71.325 189.835 72.050 ;
        RECT 190.005 71.150 190.265 71.880 ;
        RECT 190.435 71.325 190.695 72.050 ;
        RECT 190.865 71.150 191.125 71.880 ;
        RECT 191.295 71.325 191.555 72.050 ;
        RECT 191.725 71.150 191.985 71.880 ;
        RECT 192.155 71.325 192.415 72.050 ;
        RECT 192.585 71.150 192.845 72.260 ;
        RECT 193.015 71.325 193.265 72.460 ;
        RECT 193.920 72.410 195.130 72.930 ;
        RECT 193.445 71.150 193.740 72.260 ;
        RECT 195.300 72.240 196.510 72.760 ;
        RECT 193.920 71.150 196.510 72.240 ;
        RECT 196.685 72.290 196.855 72.960 ;
        RECT 197.110 72.790 197.280 72.960 ;
        RECT 197.025 72.460 197.280 72.790 ;
        RECT 197.505 72.460 197.700 72.790 ;
        RECT 196.685 71.320 197.020 72.290 ;
        RECT 197.190 71.150 197.360 72.290 ;
        RECT 197.530 71.490 197.700 72.460 ;
        RECT 197.870 71.830 198.040 72.960 ;
        RECT 198.210 72.170 198.380 72.970 ;
        RECT 198.580 72.850 198.860 73.020 ;
        RECT 198.585 72.370 198.860 72.850 ;
        RECT 199.030 72.170 199.220 73.530 ;
        RECT 199.400 73.165 199.910 73.700 ;
        RECT 200.130 72.890 200.375 73.495 ;
        RECT 200.840 73.070 201.170 73.530 ;
        RECT 201.350 73.240 201.520 73.700 ;
        RECT 201.700 73.070 202.030 73.530 ;
        RECT 202.260 73.240 202.430 73.700 ;
        RECT 202.670 73.360 203.860 73.530 ;
        RECT 202.670 73.070 203.000 73.360 ;
        RECT 203.550 73.190 203.860 73.360 ;
        RECT 204.045 73.300 204.380 73.700 ;
        RECT 200.840 72.900 203.000 73.070 ;
        RECT 199.420 72.720 200.650 72.890 ;
        RECT 198.210 72.000 199.220 72.170 ;
        RECT 199.390 72.155 200.140 72.345 ;
        RECT 197.870 71.660 198.995 71.830 ;
        RECT 199.390 71.490 199.560 72.155 ;
        RECT 200.310 71.910 200.650 72.720 ;
        RECT 200.855 72.340 201.185 72.730 ;
        RECT 201.355 72.510 202.155 72.710 ;
        RECT 202.335 72.340 202.830 72.710 ;
        RECT 200.855 72.170 202.830 72.340 ;
        RECT 203.170 72.000 203.380 73.190 ;
        RECT 204.550 73.130 204.755 73.530 ;
        RECT 204.965 73.220 205.240 73.700 ;
        RECT 205.450 73.200 205.710 73.530 ;
        RECT 203.550 72.385 203.865 73.020 ;
        RECT 204.070 72.960 204.755 73.130 ;
        RECT 197.530 71.320 199.560 71.490 ;
        RECT 199.730 71.150 199.900 71.910 ;
        RECT 200.135 71.500 200.650 71.910 ;
        RECT 200.840 71.150 201.170 72.000 ;
        RECT 201.340 71.490 201.560 72.000 ;
        RECT 201.730 71.820 203.380 72.000 ;
        RECT 201.730 71.660 202.030 71.820 ;
        RECT 202.260 71.490 202.450 71.650 ;
        RECT 201.340 71.320 202.450 71.490 ;
        RECT 202.645 71.150 202.975 71.610 ;
        RECT 203.145 71.320 203.380 71.820 ;
        RECT 203.550 71.150 203.860 72.215 ;
        RECT 204.070 71.930 204.410 72.960 ;
        RECT 204.580 72.290 204.830 72.790 ;
        RECT 205.010 72.460 205.370 73.040 ;
        RECT 205.540 72.290 205.710 73.200 ;
        RECT 205.880 72.930 209.390 73.700 ;
        RECT 209.565 72.960 209.820 73.530 ;
        RECT 209.990 73.300 210.320 73.700 ;
        RECT 210.745 73.165 211.275 73.530 ;
        RECT 210.745 73.130 210.920 73.165 ;
        RECT 209.990 72.960 210.920 73.130 ;
        RECT 205.880 72.410 207.530 72.930 ;
        RECT 204.580 72.120 205.710 72.290 ;
        RECT 207.700 72.240 209.390 72.760 ;
        RECT 204.070 71.755 204.735 71.930 ;
        RECT 204.045 71.150 204.380 71.575 ;
        RECT 204.550 71.350 204.735 71.755 ;
        RECT 204.940 71.150 205.270 71.930 ;
        RECT 205.440 71.350 205.710 72.120 ;
        RECT 205.880 71.150 209.390 72.240 ;
        RECT 209.565 72.290 209.735 72.960 ;
        RECT 209.990 72.790 210.160 72.960 ;
        RECT 209.905 72.460 210.160 72.790 ;
        RECT 210.385 72.460 210.580 72.790 ;
        RECT 209.565 71.320 209.900 72.290 ;
        RECT 210.070 71.150 210.240 72.290 ;
        RECT 210.410 71.490 210.580 72.460 ;
        RECT 210.750 71.830 210.920 72.960 ;
        RECT 211.090 72.170 211.260 72.970 ;
        RECT 211.465 72.680 211.740 73.530 ;
        RECT 211.460 72.510 211.740 72.680 ;
        RECT 211.465 72.370 211.740 72.510 ;
        RECT 211.910 72.170 212.100 73.530 ;
        RECT 212.280 73.165 212.790 73.700 ;
        RECT 213.010 72.890 213.255 73.495 ;
        RECT 213.700 72.975 213.990 73.700 ;
        RECT 214.160 72.900 214.500 73.530 ;
        RECT 214.670 72.900 214.920 73.700 ;
        RECT 215.110 73.050 215.440 73.530 ;
        RECT 215.610 73.240 215.835 73.700 ;
        RECT 216.005 73.050 216.335 73.530 ;
        RECT 212.300 72.720 213.530 72.890 ;
        RECT 211.090 72.000 212.100 72.170 ;
        RECT 212.270 72.155 213.020 72.345 ;
        RECT 210.750 71.660 211.875 71.830 ;
        RECT 212.270 71.490 212.440 72.155 ;
        RECT 213.190 71.910 213.530 72.720 ;
        RECT 214.160 72.340 214.335 72.900 ;
        RECT 215.110 72.880 216.335 73.050 ;
        RECT 216.965 72.920 217.465 73.530 ;
        RECT 217.845 73.150 218.100 73.440 ;
        RECT 218.270 73.320 218.600 73.700 ;
        RECT 217.845 72.980 218.595 73.150 ;
        RECT 214.505 72.540 215.200 72.710 ;
        RECT 210.410 71.320 212.440 71.490 ;
        RECT 212.610 71.150 212.780 71.910 ;
        RECT 213.015 71.500 213.530 71.910 ;
        RECT 213.700 71.150 213.990 72.315 ;
        RECT 214.160 72.290 214.390 72.340 ;
        RECT 215.030 72.290 215.200 72.540 ;
        RECT 215.375 72.510 215.795 72.710 ;
        RECT 215.965 72.510 216.295 72.710 ;
        RECT 216.465 72.510 216.795 72.710 ;
        RECT 216.965 72.290 217.135 72.920 ;
        RECT 217.320 72.460 217.670 72.710 ;
        RECT 214.160 71.320 214.500 72.290 ;
        RECT 214.670 71.150 214.840 72.290 ;
        RECT 215.030 72.120 217.465 72.290 ;
        RECT 217.845 72.160 218.195 72.810 ;
        RECT 215.110 71.150 215.360 71.950 ;
        RECT 216.005 71.320 216.335 72.120 ;
        RECT 216.635 71.150 216.965 71.950 ;
        RECT 217.135 71.320 217.465 72.120 ;
        RECT 218.365 71.990 218.595 72.980 ;
        RECT 217.845 71.820 218.595 71.990 ;
        RECT 217.845 71.320 218.100 71.820 ;
        RECT 218.270 71.150 218.600 71.650 ;
        RECT 218.770 71.320 218.940 73.440 ;
        RECT 219.300 73.340 219.630 73.700 ;
        RECT 219.800 73.310 220.295 73.480 ;
        RECT 220.500 73.310 221.355 73.480 ;
        RECT 219.170 72.120 219.630 73.170 ;
        RECT 219.110 71.335 219.435 72.120 ;
        RECT 219.800 71.950 219.970 73.310 ;
        RECT 220.140 72.400 220.490 73.020 ;
        RECT 220.660 72.800 221.015 73.020 ;
        RECT 220.660 72.210 220.830 72.800 ;
        RECT 221.185 72.600 221.355 73.310 ;
        RECT 222.230 73.240 222.560 73.700 ;
        RECT 222.770 73.340 223.120 73.510 ;
        RECT 221.560 72.770 222.350 73.020 ;
        RECT 222.770 72.950 223.030 73.340 ;
        RECT 223.340 73.250 224.290 73.530 ;
        RECT 224.460 73.260 224.650 73.700 ;
        RECT 224.820 73.320 225.890 73.490 ;
        RECT 222.520 72.600 222.690 72.780 ;
        RECT 219.800 71.780 220.195 71.950 ;
        RECT 220.365 71.820 220.830 72.210 ;
        RECT 221.000 72.430 222.690 72.600 ;
        RECT 220.025 71.650 220.195 71.780 ;
        RECT 221.000 71.650 221.170 72.430 ;
        RECT 222.860 72.260 223.030 72.950 ;
        RECT 221.530 72.090 223.030 72.260 ;
        RECT 223.220 72.290 223.430 73.080 ;
        RECT 223.600 72.460 223.950 73.080 ;
        RECT 224.120 72.470 224.290 73.250 ;
        RECT 224.820 73.090 224.990 73.320 ;
        RECT 224.460 72.920 224.990 73.090 ;
        RECT 224.460 72.640 224.680 72.920 ;
        RECT 225.160 72.750 225.400 73.150 ;
        RECT 224.120 72.300 224.525 72.470 ;
        RECT 224.860 72.380 225.400 72.750 ;
        RECT 225.570 72.965 225.890 73.320 ;
        RECT 226.135 73.240 226.440 73.700 ;
        RECT 226.610 72.990 226.865 73.520 ;
        RECT 225.570 72.790 225.895 72.965 ;
        RECT 225.570 72.490 226.485 72.790 ;
        RECT 225.745 72.460 226.485 72.490 ;
        RECT 223.220 72.130 223.895 72.290 ;
        RECT 224.355 72.210 224.525 72.300 ;
        RECT 223.220 72.120 224.185 72.130 ;
        RECT 222.860 71.950 223.030 72.090 ;
        RECT 219.605 71.150 219.855 71.610 ;
        RECT 220.025 71.320 220.275 71.650 ;
        RECT 220.490 71.320 221.170 71.650 ;
        RECT 221.340 71.750 222.415 71.920 ;
        RECT 222.860 71.780 223.420 71.950 ;
        RECT 223.725 71.830 224.185 72.120 ;
        RECT 224.355 72.040 225.575 72.210 ;
        RECT 221.340 71.410 221.510 71.750 ;
        RECT 221.745 71.150 222.075 71.580 ;
        RECT 222.245 71.410 222.415 71.750 ;
        RECT 222.710 71.150 223.080 71.610 ;
        RECT 223.250 71.320 223.420 71.780 ;
        RECT 224.355 71.660 224.525 72.040 ;
        RECT 225.745 71.870 225.915 72.460 ;
        RECT 226.655 72.340 226.865 72.990 ;
        RECT 227.040 72.930 229.630 73.700 ;
        RECT 229.805 72.935 230.260 73.700 ;
        RECT 230.535 73.320 231.835 73.530 ;
        RECT 232.090 73.340 232.420 73.700 ;
        RECT 231.665 73.170 231.835 73.320 ;
        RECT 232.590 73.200 232.850 73.530 ;
        RECT 227.040 72.410 228.250 72.930 ;
        RECT 223.655 71.320 224.525 71.660 ;
        RECT 225.115 71.700 225.915 71.870 ;
        RECT 224.695 71.150 224.945 71.610 ;
        RECT 225.115 71.410 225.285 71.700 ;
        RECT 225.465 71.150 225.795 71.530 ;
        RECT 226.135 71.150 226.440 72.290 ;
        RECT 226.610 71.460 226.865 72.340 ;
        RECT 228.420 72.240 229.630 72.760 ;
        RECT 230.735 72.710 230.955 73.110 ;
        RECT 229.800 72.510 230.290 72.710 ;
        RECT 230.480 72.500 230.955 72.710 ;
        RECT 231.200 72.710 231.410 73.110 ;
        RECT 231.665 73.045 232.420 73.170 ;
        RECT 231.665 73.000 232.510 73.045 ;
        RECT 232.240 72.880 232.510 73.000 ;
        RECT 231.200 72.500 231.530 72.710 ;
        RECT 231.700 72.440 232.110 72.745 ;
        RECT 227.040 71.150 229.630 72.240 ;
        RECT 229.805 72.270 230.980 72.330 ;
        RECT 232.340 72.305 232.510 72.880 ;
        RECT 232.310 72.270 232.510 72.305 ;
        RECT 229.805 72.160 232.510 72.270 ;
        RECT 229.805 71.540 230.060 72.160 ;
        RECT 230.650 72.100 232.450 72.160 ;
        RECT 230.650 72.070 230.980 72.100 ;
        RECT 232.680 72.000 232.850 73.200 ;
        RECT 233.020 73.155 238.365 73.700 ;
        RECT 234.605 72.325 234.945 73.155 ;
        RECT 239.460 72.975 239.750 73.700 ;
        RECT 240.010 73.050 240.180 73.530 ;
        RECT 240.350 73.220 240.680 73.700 ;
        RECT 240.905 73.280 242.440 73.530 ;
        RECT 240.905 73.050 241.075 73.280 ;
        RECT 240.010 72.880 241.075 73.050 ;
        RECT 230.310 71.900 230.495 71.990 ;
        RECT 231.085 71.900 231.920 71.910 ;
        RECT 230.310 71.700 231.920 71.900 ;
        RECT 230.310 71.660 230.540 71.700 ;
        RECT 229.805 71.320 230.140 71.540 ;
        RECT 231.145 71.150 231.500 71.530 ;
        RECT 231.670 71.320 231.920 71.700 ;
        RECT 232.170 71.150 232.420 71.930 ;
        RECT 232.590 71.320 232.850 72.000 ;
        RECT 236.425 71.585 236.775 72.835 ;
        RECT 241.255 72.710 241.535 73.110 ;
        RECT 239.925 72.500 240.275 72.710 ;
        RECT 240.445 72.510 240.890 72.710 ;
        RECT 241.060 72.510 241.535 72.710 ;
        RECT 241.805 72.710 242.090 73.110 ;
        RECT 242.270 73.050 242.440 73.280 ;
        RECT 242.610 73.220 242.940 73.700 ;
        RECT 243.155 73.200 243.410 73.530 ;
        RECT 243.225 73.120 243.410 73.200 ;
        RECT 242.270 72.880 243.070 73.050 ;
        RECT 241.805 72.510 242.135 72.710 ;
        RECT 242.305 72.680 242.670 72.710 ;
        RECT 242.305 72.510 242.680 72.680 ;
        RECT 242.900 72.330 243.070 72.880 ;
        RECT 233.020 71.150 238.365 71.585 ;
        RECT 239.460 71.150 239.750 72.315 ;
        RECT 240.010 72.160 243.070 72.330 ;
        RECT 240.010 71.320 240.180 72.160 ;
        RECT 243.240 71.990 243.410 73.120 ;
        RECT 240.350 71.490 240.680 71.990 ;
        RECT 240.850 71.750 242.485 71.990 ;
        RECT 240.850 71.660 241.080 71.750 ;
        RECT 241.190 71.490 241.520 71.530 ;
        RECT 240.350 71.320 241.520 71.490 ;
        RECT 241.710 71.150 242.065 71.570 ;
        RECT 242.235 71.320 242.485 71.750 ;
        RECT 242.655 71.150 242.985 71.910 ;
        RECT 243.155 71.320 243.410 71.990 ;
        RECT 243.620 73.200 243.875 73.530 ;
        RECT 244.090 73.220 244.420 73.700 ;
        RECT 244.590 73.280 246.125 73.530 ;
        RECT 243.620 73.120 243.805 73.200 ;
        RECT 243.620 72.000 243.790 73.120 ;
        RECT 244.590 73.050 244.760 73.280 ;
        RECT 243.960 72.880 244.760 73.050 ;
        RECT 243.960 72.330 244.130 72.880 ;
        RECT 244.940 72.710 245.225 73.110 ;
        RECT 244.360 72.680 244.725 72.710 ;
        RECT 244.350 72.510 244.725 72.680 ;
        RECT 244.895 72.510 245.225 72.710 ;
        RECT 245.495 72.710 245.775 73.110 ;
        RECT 245.955 73.050 246.125 73.280 ;
        RECT 246.350 73.220 246.680 73.700 ;
        RECT 246.850 73.050 247.020 73.530 ;
        RECT 247.280 73.155 252.625 73.700 ;
        RECT 245.955 72.880 247.020 73.050 ;
        RECT 245.495 72.510 245.970 72.710 ;
        RECT 246.140 72.510 246.585 72.710 ;
        RECT 246.755 72.500 247.105 72.710 ;
        RECT 243.960 72.160 247.020 72.330 ;
        RECT 248.865 72.325 249.205 73.155 ;
        RECT 252.800 72.930 256.310 73.700 ;
        RECT 256.485 72.935 256.940 73.700 ;
        RECT 257.215 73.320 258.515 73.530 ;
        RECT 258.770 73.340 259.100 73.700 ;
        RECT 258.345 73.170 258.515 73.320 ;
        RECT 259.270 73.200 259.530 73.530 ;
        RECT 243.620 71.990 243.830 72.000 ;
        RECT 243.620 71.320 243.875 71.990 ;
        RECT 244.045 71.150 244.375 71.910 ;
        RECT 244.545 71.750 246.180 71.990 ;
        RECT 244.545 71.320 244.795 71.750 ;
        RECT 245.950 71.660 246.180 71.750 ;
        RECT 244.965 71.150 245.320 71.570 ;
        RECT 245.510 71.490 245.840 71.530 ;
        RECT 246.350 71.490 246.680 71.990 ;
        RECT 245.510 71.320 246.680 71.490 ;
        RECT 246.850 71.320 247.020 72.160 ;
        RECT 250.685 71.585 251.035 72.835 ;
        RECT 252.800 72.410 254.450 72.930 ;
        RECT 254.620 72.240 256.310 72.760 ;
        RECT 257.415 72.710 257.635 73.110 ;
        RECT 256.480 72.510 256.970 72.710 ;
        RECT 257.160 72.500 257.635 72.710 ;
        RECT 257.880 72.710 258.090 73.110 ;
        RECT 258.345 73.045 259.100 73.170 ;
        RECT 258.345 73.000 259.190 73.045 ;
        RECT 258.920 72.880 259.190 73.000 ;
        RECT 257.880 72.500 258.210 72.710 ;
        RECT 258.380 72.440 258.790 72.745 ;
        RECT 247.280 71.150 252.625 71.585 ;
        RECT 252.800 71.150 256.310 72.240 ;
        RECT 256.485 72.270 257.660 72.330 ;
        RECT 259.020 72.305 259.190 72.880 ;
        RECT 258.990 72.270 259.190 72.305 ;
        RECT 256.485 72.160 259.190 72.270 ;
        RECT 256.485 71.540 256.740 72.160 ;
        RECT 257.330 72.100 259.130 72.160 ;
        RECT 257.330 72.070 257.660 72.100 ;
        RECT 259.360 72.000 259.530 73.200 ;
        RECT 259.790 73.050 259.960 73.530 ;
        RECT 260.130 73.220 260.460 73.700 ;
        RECT 260.685 73.280 262.220 73.530 ;
        RECT 260.685 73.050 260.855 73.280 ;
        RECT 259.790 72.880 260.855 73.050 ;
        RECT 261.035 72.710 261.315 73.110 ;
        RECT 259.705 72.500 260.055 72.710 ;
        RECT 260.225 72.510 260.670 72.710 ;
        RECT 260.840 72.510 261.315 72.710 ;
        RECT 261.585 72.710 261.870 73.110 ;
        RECT 262.050 73.050 262.220 73.280 ;
        RECT 262.390 73.220 262.720 73.700 ;
        RECT 262.935 73.200 263.190 73.530 ;
        RECT 263.005 73.120 263.190 73.200 ;
        RECT 262.050 72.880 262.850 73.050 ;
        RECT 261.585 72.510 261.915 72.710 ;
        RECT 262.085 72.510 262.450 72.710 ;
        RECT 262.680 72.330 262.850 72.880 ;
        RECT 256.990 71.900 257.175 71.990 ;
        RECT 257.765 71.900 258.600 71.910 ;
        RECT 256.990 71.700 258.600 71.900 ;
        RECT 256.990 71.660 257.220 71.700 ;
        RECT 256.485 71.320 256.820 71.540 ;
        RECT 257.825 71.150 258.180 71.530 ;
        RECT 258.350 71.320 258.600 71.700 ;
        RECT 258.850 71.150 259.100 71.930 ;
        RECT 259.270 71.320 259.530 72.000 ;
        RECT 259.790 72.160 262.850 72.330 ;
        RECT 259.790 71.320 259.960 72.160 ;
        RECT 263.020 72.000 263.190 73.120 ;
        RECT 263.380 72.930 265.050 73.700 ;
        RECT 265.220 72.975 265.510 73.700 ;
        RECT 265.680 73.200 265.940 73.530 ;
        RECT 266.110 73.340 266.440 73.700 ;
        RECT 266.695 73.320 267.995 73.530 ;
        RECT 263.380 72.410 264.130 72.930 ;
        RECT 264.300 72.240 265.050 72.760 ;
        RECT 262.980 71.990 263.190 72.000 ;
        RECT 260.130 71.490 260.460 71.990 ;
        RECT 260.630 71.750 262.265 71.990 ;
        RECT 260.630 71.660 260.860 71.750 ;
        RECT 260.970 71.490 261.300 71.530 ;
        RECT 260.130 71.320 261.300 71.490 ;
        RECT 261.490 71.150 261.845 71.570 ;
        RECT 262.015 71.320 262.265 71.750 ;
        RECT 262.435 71.150 262.765 71.910 ;
        RECT 262.935 71.320 263.190 71.990 ;
        RECT 263.380 71.150 265.050 72.240 ;
        RECT 265.220 71.150 265.510 72.315 ;
        RECT 265.680 72.000 265.850 73.200 ;
        RECT 266.695 73.170 266.865 73.320 ;
        RECT 266.110 73.045 266.865 73.170 ;
        RECT 266.020 73.000 266.865 73.045 ;
        RECT 266.020 72.880 266.290 73.000 ;
        RECT 266.020 72.305 266.190 72.880 ;
        RECT 266.420 72.440 266.830 72.745 ;
        RECT 267.120 72.710 267.330 73.110 ;
        RECT 267.000 72.500 267.330 72.710 ;
        RECT 267.575 72.710 267.795 73.110 ;
        RECT 268.270 72.935 268.725 73.700 ;
        RECT 268.900 73.155 274.245 73.700 ;
        RECT 267.575 72.500 268.050 72.710 ;
        RECT 268.240 72.510 268.730 72.710 ;
        RECT 266.020 72.270 266.220 72.305 ;
        RECT 267.550 72.270 268.725 72.330 ;
        RECT 270.485 72.325 270.825 73.155 ;
        RECT 274.420 72.950 275.630 73.700 ;
        RECT 275.800 73.070 276.140 73.530 ;
        RECT 276.310 73.240 276.480 73.700 ;
        RECT 277.110 73.265 277.470 73.530 ;
        RECT 277.115 73.260 277.470 73.265 ;
        RECT 277.120 73.250 277.470 73.260 ;
        RECT 277.125 73.245 277.470 73.250 ;
        RECT 277.130 73.235 277.470 73.245 ;
        RECT 277.710 73.240 277.880 73.700 ;
        RECT 277.135 73.230 277.470 73.235 ;
        RECT 277.145 73.220 277.470 73.230 ;
        RECT 277.155 73.210 277.470 73.220 ;
        RECT 276.650 73.070 276.980 73.150 ;
        RECT 266.020 72.160 268.725 72.270 ;
        RECT 266.080 72.100 267.880 72.160 ;
        RECT 267.550 72.070 267.880 72.100 ;
        RECT 265.680 71.320 265.940 72.000 ;
        RECT 266.110 71.150 266.360 71.930 ;
        RECT 266.610 71.900 267.445 71.910 ;
        RECT 268.035 71.900 268.220 71.990 ;
        RECT 266.610 71.700 268.220 71.900 ;
        RECT 266.610 71.320 266.860 71.700 ;
        RECT 267.990 71.660 268.220 71.700 ;
        RECT 268.470 71.540 268.725 72.160 ;
        RECT 272.305 71.585 272.655 72.835 ;
        RECT 274.420 72.410 274.940 72.950 ;
        RECT 275.800 72.880 276.980 73.070 ;
        RECT 277.170 73.070 277.470 73.210 ;
        RECT 277.170 72.880 277.880 73.070 ;
        RECT 275.110 72.240 275.630 72.780 ;
        RECT 267.030 71.150 267.385 71.530 ;
        RECT 268.390 71.320 268.725 71.540 ;
        RECT 268.900 71.150 274.245 71.585 ;
        RECT 274.420 71.150 275.630 72.240 ;
        RECT 275.800 72.510 276.130 72.710 ;
        RECT 276.440 72.690 276.770 72.710 ;
        RECT 276.320 72.510 276.770 72.690 ;
        RECT 275.800 72.170 276.030 72.510 ;
        RECT 275.810 71.150 276.140 71.870 ;
        RECT 276.320 71.395 276.535 72.510 ;
        RECT 276.940 72.480 277.410 72.710 ;
        RECT 277.595 72.310 277.880 72.880 ;
        RECT 278.050 72.755 278.390 73.530 ;
        RECT 278.565 73.150 278.820 73.440 ;
        RECT 278.990 73.320 279.320 73.700 ;
        RECT 278.565 72.980 279.315 73.150 ;
        RECT 276.730 72.095 277.880 72.310 ;
        RECT 276.730 71.320 277.060 72.095 ;
        RECT 277.230 71.150 277.940 71.925 ;
        RECT 278.110 71.320 278.390 72.755 ;
        RECT 278.565 72.160 278.915 72.810 ;
        RECT 279.085 71.990 279.315 72.980 ;
        RECT 278.565 71.820 279.315 71.990 ;
        RECT 278.565 71.320 278.820 71.820 ;
        RECT 278.990 71.150 279.320 71.650 ;
        RECT 279.490 71.320 279.660 73.440 ;
        RECT 280.020 73.340 280.350 73.700 ;
        RECT 280.520 73.310 281.015 73.480 ;
        RECT 281.220 73.310 282.075 73.480 ;
        RECT 279.890 72.120 280.350 73.170 ;
        RECT 279.830 71.335 280.155 72.120 ;
        RECT 280.520 71.950 280.690 73.310 ;
        RECT 280.860 72.400 281.210 73.020 ;
        RECT 281.380 72.800 281.735 73.020 ;
        RECT 281.380 72.210 281.550 72.800 ;
        RECT 281.905 72.600 282.075 73.310 ;
        RECT 282.950 73.240 283.280 73.700 ;
        RECT 283.490 73.340 283.840 73.510 ;
        RECT 282.280 72.770 283.070 73.020 ;
        RECT 283.490 72.950 283.750 73.340 ;
        RECT 284.060 73.250 285.010 73.530 ;
        RECT 285.180 73.260 285.370 73.700 ;
        RECT 285.540 73.320 286.610 73.490 ;
        RECT 283.240 72.600 283.410 72.780 ;
        RECT 280.520 71.780 280.915 71.950 ;
        RECT 281.085 71.820 281.550 72.210 ;
        RECT 281.720 72.430 283.410 72.600 ;
        RECT 280.745 71.650 280.915 71.780 ;
        RECT 281.720 71.650 281.890 72.430 ;
        RECT 283.580 72.260 283.750 72.950 ;
        RECT 282.250 72.090 283.750 72.260 ;
        RECT 283.940 72.290 284.150 73.080 ;
        RECT 284.320 72.460 284.670 73.080 ;
        RECT 284.840 72.470 285.010 73.250 ;
        RECT 285.540 73.090 285.710 73.320 ;
        RECT 285.180 72.920 285.710 73.090 ;
        RECT 285.180 72.640 285.400 72.920 ;
        RECT 285.880 72.750 286.120 73.150 ;
        RECT 284.840 72.300 285.245 72.470 ;
        RECT 285.580 72.380 286.120 72.750 ;
        RECT 286.290 72.965 286.610 73.320 ;
        RECT 286.855 73.240 287.160 73.700 ;
        RECT 287.330 72.990 287.585 73.520 ;
        RECT 288.890 73.010 289.220 73.700 ;
        RECT 289.680 73.105 290.300 73.530 ;
        RECT 290.470 73.210 290.800 73.700 ;
        RECT 286.290 72.790 286.615 72.965 ;
        RECT 286.290 72.490 287.205 72.790 ;
        RECT 286.465 72.460 287.205 72.490 ;
        RECT 283.940 72.130 284.615 72.290 ;
        RECT 285.075 72.210 285.245 72.300 ;
        RECT 283.940 72.120 284.905 72.130 ;
        RECT 283.580 71.950 283.750 72.090 ;
        RECT 280.325 71.150 280.575 71.610 ;
        RECT 280.745 71.320 280.995 71.650 ;
        RECT 281.210 71.320 281.890 71.650 ;
        RECT 282.060 71.750 283.135 71.920 ;
        RECT 283.580 71.780 284.140 71.950 ;
        RECT 284.445 71.830 284.905 72.120 ;
        RECT 285.075 72.040 286.295 72.210 ;
        RECT 282.060 71.410 282.230 71.750 ;
        RECT 282.465 71.150 282.795 71.580 ;
        RECT 282.965 71.410 283.135 71.750 ;
        RECT 283.430 71.150 283.800 71.610 ;
        RECT 283.970 71.320 284.140 71.780 ;
        RECT 285.075 71.660 285.245 72.040 ;
        RECT 286.465 71.870 286.635 72.460 ;
        RECT 287.375 72.340 287.585 72.990 ;
        RECT 289.940 72.770 290.300 73.105 ;
        RECT 284.375 71.320 285.245 71.660 ;
        RECT 285.835 71.700 286.635 71.870 ;
        RECT 285.415 71.150 285.665 71.610 ;
        RECT 285.835 71.410 286.005 71.700 ;
        RECT 286.185 71.150 286.515 71.530 ;
        RECT 286.855 71.150 287.160 72.290 ;
        RECT 287.330 71.460 287.585 72.340 ;
        RECT 288.880 72.490 290.300 72.770 ;
        RECT 288.350 71.150 288.680 72.320 ;
        RECT 288.880 71.320 289.210 72.490 ;
        RECT 289.410 71.150 289.740 72.320 ;
        RECT 289.940 71.320 290.300 72.490 ;
        RECT 290.470 72.460 290.810 73.040 ;
        RECT 290.980 72.975 291.270 73.700 ;
        RECT 291.440 72.930 293.110 73.700 ;
        RECT 293.285 72.990 293.540 73.520 ;
        RECT 293.710 73.240 294.015 73.700 ;
        RECT 294.260 73.320 295.330 73.490 ;
        RECT 291.440 72.410 292.190 72.930 ;
        RECT 290.470 71.150 290.800 72.290 ;
        RECT 290.980 71.150 291.270 72.315 ;
        RECT 292.360 72.240 293.110 72.760 ;
        RECT 291.440 71.150 293.110 72.240 ;
        RECT 293.285 72.340 293.495 72.990 ;
        RECT 294.260 72.965 294.580 73.320 ;
        RECT 294.255 72.790 294.580 72.965 ;
        RECT 293.665 72.490 294.580 72.790 ;
        RECT 294.750 72.750 294.990 73.150 ;
        RECT 295.160 73.090 295.330 73.320 ;
        RECT 295.500 73.260 295.690 73.700 ;
        RECT 295.860 73.250 296.810 73.530 ;
        RECT 297.030 73.340 297.380 73.510 ;
        RECT 295.160 72.920 295.690 73.090 ;
        RECT 293.665 72.460 294.405 72.490 ;
        RECT 293.285 71.460 293.540 72.340 ;
        RECT 293.710 71.150 294.015 72.290 ;
        RECT 294.235 71.870 294.405 72.460 ;
        RECT 294.750 72.380 295.290 72.750 ;
        RECT 295.470 72.640 295.690 72.920 ;
        RECT 295.860 72.470 296.030 73.250 ;
        RECT 295.625 72.300 296.030 72.470 ;
        RECT 296.200 72.460 296.550 73.080 ;
        RECT 295.625 72.210 295.795 72.300 ;
        RECT 296.720 72.290 296.930 73.080 ;
        RECT 294.575 72.040 295.795 72.210 ;
        RECT 296.255 72.130 296.930 72.290 ;
        RECT 294.235 71.700 295.035 71.870 ;
        RECT 294.355 71.150 294.685 71.530 ;
        RECT 294.865 71.410 295.035 71.700 ;
        RECT 295.625 71.660 295.795 72.040 ;
        RECT 295.965 72.120 296.930 72.130 ;
        RECT 297.120 72.950 297.380 73.340 ;
        RECT 297.590 73.240 297.920 73.700 ;
        RECT 298.795 73.310 299.650 73.480 ;
        RECT 299.855 73.310 300.350 73.480 ;
        RECT 300.520 73.340 300.850 73.700 ;
        RECT 297.120 72.260 297.290 72.950 ;
        RECT 297.460 72.600 297.630 72.780 ;
        RECT 297.800 72.770 298.590 73.020 ;
        RECT 298.795 72.600 298.965 73.310 ;
        RECT 299.135 72.800 299.490 73.020 ;
        RECT 297.460 72.430 299.150 72.600 ;
        RECT 295.965 71.830 296.425 72.120 ;
        RECT 297.120 72.090 298.620 72.260 ;
        RECT 297.120 71.950 297.290 72.090 ;
        RECT 296.730 71.780 297.290 71.950 ;
        RECT 295.205 71.150 295.455 71.610 ;
        RECT 295.625 71.320 296.495 71.660 ;
        RECT 296.730 71.320 296.900 71.780 ;
        RECT 297.735 71.750 298.810 71.920 ;
        RECT 297.070 71.150 297.440 71.610 ;
        RECT 297.735 71.410 297.905 71.750 ;
        RECT 298.075 71.150 298.405 71.580 ;
        RECT 298.640 71.410 298.810 71.750 ;
        RECT 298.980 71.650 299.150 72.430 ;
        RECT 299.320 72.210 299.490 72.800 ;
        RECT 299.660 72.400 300.010 73.020 ;
        RECT 299.320 71.820 299.785 72.210 ;
        RECT 300.180 71.950 300.350 73.310 ;
        RECT 300.520 72.120 300.980 73.170 ;
        RECT 299.955 71.780 300.350 71.950 ;
        RECT 299.955 71.650 300.125 71.780 ;
        RECT 298.980 71.320 299.660 71.650 ;
        RECT 299.875 71.320 300.125 71.650 ;
        RECT 300.295 71.150 300.545 71.610 ;
        RECT 300.715 71.335 301.040 72.120 ;
        RECT 301.210 71.320 301.380 73.440 ;
        RECT 301.550 73.320 301.880 73.700 ;
        RECT 302.050 73.150 302.305 73.440 ;
        RECT 301.555 72.980 302.305 73.150 ;
        RECT 301.555 71.990 301.785 72.980 ;
        RECT 302.485 72.960 302.740 73.530 ;
        RECT 302.910 73.300 303.240 73.700 ;
        RECT 303.665 73.165 304.195 73.530 ;
        RECT 304.385 73.360 304.660 73.530 ;
        RECT 304.380 73.190 304.660 73.360 ;
        RECT 303.665 73.130 303.840 73.165 ;
        RECT 302.910 72.960 303.840 73.130 ;
        RECT 301.955 72.160 302.305 72.810 ;
        RECT 302.485 72.290 302.655 72.960 ;
        RECT 302.910 72.790 303.080 72.960 ;
        RECT 302.825 72.460 303.080 72.790 ;
        RECT 303.305 72.460 303.500 72.790 ;
        RECT 301.555 71.820 302.305 71.990 ;
        RECT 301.550 71.150 301.880 71.650 ;
        RECT 302.050 71.320 302.305 71.820 ;
        RECT 302.485 71.320 302.820 72.290 ;
        RECT 302.990 71.150 303.160 72.290 ;
        RECT 303.330 71.490 303.500 72.460 ;
        RECT 303.670 71.830 303.840 72.960 ;
        RECT 304.010 72.170 304.180 72.970 ;
        RECT 304.385 72.370 304.660 73.190 ;
        RECT 304.830 72.170 305.020 73.530 ;
        RECT 305.200 73.165 305.710 73.700 ;
        RECT 305.930 72.890 306.175 73.495 ;
        RECT 305.220 72.720 306.450 72.890 ;
        RECT 306.625 72.860 306.885 73.700 ;
        RECT 307.060 72.955 307.315 73.530 ;
        RECT 307.485 73.320 307.815 73.700 ;
        RECT 308.030 73.150 308.200 73.530 ;
        RECT 307.485 72.980 308.200 73.150 ;
        RECT 304.010 72.000 305.020 72.170 ;
        RECT 305.190 72.155 305.940 72.345 ;
        RECT 303.670 71.660 304.795 71.830 ;
        RECT 305.190 71.490 305.360 72.155 ;
        RECT 306.110 71.910 306.450 72.720 ;
        RECT 303.330 71.320 305.360 71.490 ;
        RECT 305.530 71.150 305.700 71.910 ;
        RECT 305.935 71.500 306.450 71.910 ;
        RECT 306.625 71.150 306.885 72.300 ;
        RECT 307.060 72.225 307.230 72.955 ;
        RECT 307.485 72.790 307.655 72.980 ;
        RECT 308.460 72.950 309.670 73.700 ;
        RECT 309.840 72.950 311.050 73.700 ;
        RECT 307.400 72.460 307.655 72.790 ;
        RECT 307.485 72.250 307.655 72.460 ;
        RECT 307.935 72.430 308.290 72.800 ;
        RECT 308.460 72.410 308.980 72.950 ;
        RECT 307.060 71.320 307.315 72.225 ;
        RECT 307.485 72.080 308.200 72.250 ;
        RECT 309.150 72.240 309.670 72.780 ;
        RECT 307.485 71.150 307.815 71.910 ;
        RECT 308.030 71.320 308.200 72.080 ;
        RECT 308.460 71.150 309.670 72.240 ;
        RECT 309.840 72.240 310.360 72.780 ;
        RECT 310.530 72.410 311.050 72.950 ;
        RECT 309.840 71.150 311.050 72.240 ;
        RECT 162.095 70.980 311.135 71.150 ;
        RECT 162.180 69.890 163.390 70.980 ;
        RECT 163.560 70.545 168.905 70.980 ;
        RECT 162.180 69.180 162.700 69.720 ;
        RECT 162.870 69.350 163.390 69.890 ;
        RECT 162.180 68.430 163.390 69.180 ;
        RECT 165.145 68.975 165.485 69.805 ;
        RECT 166.965 69.295 167.315 70.545 ;
        RECT 169.080 69.890 170.750 70.980 ;
        RECT 169.080 69.200 169.830 69.720 ;
        RECT 170.000 69.370 170.750 69.890 ;
        RECT 170.925 69.840 171.260 70.810 ;
        RECT 171.430 69.840 171.600 70.980 ;
        RECT 171.770 70.640 173.800 70.810 ;
        RECT 163.560 68.430 168.905 68.975 ;
        RECT 169.080 68.430 170.750 69.200 ;
        RECT 170.925 69.170 171.095 69.840 ;
        RECT 171.770 69.670 171.940 70.640 ;
        RECT 171.265 69.340 171.520 69.670 ;
        RECT 171.745 69.340 171.940 69.670 ;
        RECT 172.110 70.300 173.235 70.470 ;
        RECT 171.350 69.170 171.520 69.340 ;
        RECT 172.110 69.170 172.280 70.300 ;
        RECT 170.925 68.600 171.180 69.170 ;
        RECT 171.350 69.000 172.280 69.170 ;
        RECT 172.450 69.960 173.460 70.130 ;
        RECT 172.450 69.160 172.620 69.960 ;
        RECT 172.105 68.965 172.280 69.000 ;
        RECT 171.350 68.430 171.680 68.830 ;
        RECT 172.105 68.600 172.635 68.965 ;
        RECT 172.825 68.940 173.100 69.760 ;
        RECT 172.820 68.770 173.100 68.940 ;
        RECT 172.825 68.600 173.100 68.770 ;
        RECT 173.270 68.600 173.460 69.960 ;
        RECT 173.630 69.975 173.800 70.640 ;
        RECT 173.970 70.220 174.140 70.980 ;
        RECT 174.375 70.220 174.890 70.630 ;
        RECT 173.630 69.785 174.380 69.975 ;
        RECT 174.550 69.410 174.890 70.220 ;
        RECT 175.060 69.815 175.350 70.980 ;
        RECT 175.525 69.840 175.860 70.810 ;
        RECT 176.030 69.840 176.200 70.980 ;
        RECT 176.370 70.640 178.400 70.810 ;
        RECT 173.660 69.240 174.890 69.410 ;
        RECT 173.640 68.430 174.150 68.965 ;
        RECT 174.370 68.635 174.615 69.240 ;
        RECT 175.525 69.170 175.695 69.840 ;
        RECT 176.370 69.670 176.540 70.640 ;
        RECT 175.865 69.340 176.120 69.670 ;
        RECT 176.345 69.340 176.540 69.670 ;
        RECT 176.710 70.300 177.835 70.470 ;
        RECT 175.950 69.170 176.120 69.340 ;
        RECT 176.710 69.170 176.880 70.300 ;
        RECT 175.060 68.430 175.350 69.155 ;
        RECT 175.525 68.600 175.780 69.170 ;
        RECT 175.950 69.000 176.880 69.170 ;
        RECT 177.050 69.960 178.060 70.130 ;
        RECT 177.050 69.160 177.220 69.960 ;
        RECT 176.705 68.965 176.880 69.000 ;
        RECT 175.950 68.430 176.280 68.830 ;
        RECT 176.705 68.600 177.235 68.965 ;
        RECT 177.425 68.940 177.700 69.760 ;
        RECT 177.420 68.770 177.700 68.940 ;
        RECT 177.425 68.600 177.700 68.770 ;
        RECT 177.870 68.600 178.060 69.960 ;
        RECT 178.230 69.975 178.400 70.640 ;
        RECT 178.570 70.220 178.740 70.980 ;
        RECT 178.975 70.220 179.490 70.630 ;
        RECT 178.230 69.785 178.980 69.975 ;
        RECT 179.150 69.410 179.490 70.220 ;
        RECT 179.660 69.890 183.170 70.980 ;
        RECT 183.805 70.180 184.120 70.980 ;
        RECT 184.385 70.625 185.465 70.795 ;
        RECT 184.385 70.010 184.555 70.625 ;
        RECT 178.260 69.240 179.490 69.410 ;
        RECT 178.240 68.430 178.750 68.965 ;
        RECT 178.970 68.635 179.215 69.240 ;
        RECT 179.660 69.200 181.310 69.720 ;
        RECT 181.480 69.370 183.170 69.890 ;
        RECT 179.660 68.430 183.170 69.200 ;
        RECT 183.800 69.000 184.070 70.010 ;
        RECT 184.240 69.840 184.555 70.010 ;
        RECT 184.240 69.170 184.410 69.840 ;
        RECT 184.725 69.670 184.960 70.350 ;
        RECT 185.130 69.840 185.465 70.625 ;
        RECT 186.370 70.470 186.700 70.980 ;
        RECT 185.640 70.130 187.600 70.300 ;
        RECT 184.580 69.340 184.960 69.670 ;
        RECT 185.130 69.340 185.465 69.670 ;
        RECT 185.640 69.170 185.810 70.130 ;
        RECT 185.980 69.340 186.330 69.960 ;
        RECT 186.500 69.340 186.840 69.960 ;
        RECT 187.010 69.340 187.250 69.960 ;
        RECT 187.430 69.590 187.600 70.130 ;
        RECT 187.770 69.790 188.230 70.800 ;
        RECT 187.430 69.420 187.890 69.590 ;
        RECT 188.060 69.170 188.230 69.790 ;
        RECT 184.240 69.000 185.465 69.170 ;
        RECT 185.640 69.000 186.135 69.170 ;
        RECT 183.870 68.430 184.200 68.830 ;
        RECT 184.370 68.730 184.540 69.000 ;
        RECT 184.710 68.430 185.040 68.830 ;
        RECT 185.210 68.730 185.465 69.000 ;
        RECT 185.965 68.750 186.135 69.000 ;
        RECT 186.370 68.430 186.700 69.170 ;
        RECT 186.870 69.000 188.230 69.170 ;
        RECT 186.870 68.655 187.040 69.000 ;
        RECT 187.210 68.430 187.540 68.830 ;
        RECT 187.710 68.600 188.230 69.000 ;
        RECT 188.405 69.840 188.740 70.810 ;
        RECT 188.910 69.840 189.080 70.980 ;
        RECT 189.250 70.640 191.280 70.810 ;
        RECT 188.405 69.170 188.575 69.840 ;
        RECT 189.250 69.670 189.420 70.640 ;
        RECT 188.745 69.340 189.000 69.670 ;
        RECT 189.225 69.340 189.420 69.670 ;
        RECT 189.590 70.300 190.715 70.470 ;
        RECT 188.830 69.170 189.000 69.340 ;
        RECT 189.590 69.170 189.760 70.300 ;
        RECT 188.405 68.600 188.660 69.170 ;
        RECT 188.830 69.000 189.760 69.170 ;
        RECT 189.930 69.960 190.940 70.130 ;
        RECT 189.930 69.160 190.100 69.960 ;
        RECT 189.585 68.965 189.760 69.000 ;
        RECT 188.830 68.430 189.160 68.830 ;
        RECT 189.585 68.600 190.115 68.965 ;
        RECT 190.305 68.940 190.580 69.760 ;
        RECT 190.300 68.770 190.580 68.940 ;
        RECT 190.305 68.600 190.580 68.770 ;
        RECT 190.750 68.600 190.940 69.960 ;
        RECT 191.110 69.975 191.280 70.640 ;
        RECT 191.450 70.220 191.620 70.980 ;
        RECT 191.855 70.220 192.370 70.630 ;
        RECT 191.110 69.785 191.860 69.975 ;
        RECT 192.030 69.410 192.370 70.220 ;
        RECT 193.510 69.885 193.760 70.980 ;
        RECT 194.495 70.640 196.560 70.810 ;
        RECT 193.930 69.800 194.285 70.215 ;
        RECT 194.495 69.800 194.740 70.640 ;
        RECT 194.115 69.630 194.285 69.800 ;
        RECT 193.460 69.420 193.945 69.630 ;
        RECT 194.115 69.420 194.740 69.630 ;
        RECT 191.140 69.240 192.370 69.410 ;
        RECT 194.115 69.250 194.285 69.420 ;
        RECT 194.910 69.250 195.160 70.470 ;
        RECT 195.330 69.800 195.600 70.640 ;
        RECT 195.890 69.970 196.140 70.470 ;
        RECT 196.310 70.140 196.560 70.640 ;
        RECT 196.730 69.970 196.980 70.810 ;
        RECT 197.150 70.140 197.400 70.980 ;
        RECT 197.570 69.970 197.885 70.810 ;
        RECT 195.890 69.800 197.885 69.970 ;
        RECT 198.060 69.890 200.650 70.980 ;
        RECT 195.335 69.420 196.840 69.630 ;
        RECT 197.010 69.420 197.865 69.630 ;
        RECT 191.120 68.430 191.630 68.965 ;
        RECT 191.850 68.635 192.095 69.240 ;
        RECT 193.470 68.430 193.760 69.170 ;
        RECT 193.930 68.725 194.285 69.250 ;
        RECT 194.495 68.430 194.700 69.240 ;
        RECT 194.870 69.070 197.440 69.250 ;
        RECT 194.870 68.600 195.200 69.070 ;
        RECT 195.370 68.430 196.100 68.900 ;
        RECT 196.270 68.600 196.600 69.070 ;
        RECT 196.770 68.430 196.940 68.900 ;
        RECT 197.110 68.600 197.440 69.070 ;
        RECT 197.610 68.430 197.885 69.250 ;
        RECT 198.060 69.200 199.270 69.720 ;
        RECT 199.440 69.370 200.650 69.890 ;
        RECT 200.820 69.815 201.110 70.980 ;
        RECT 201.280 70.545 206.625 70.980 ;
        RECT 198.060 68.430 200.650 69.200 ;
        RECT 200.820 68.430 201.110 69.155 ;
        RECT 202.865 68.975 203.205 69.805 ;
        RECT 204.685 69.295 205.035 70.545 ;
        RECT 207.265 70.310 207.520 70.810 ;
        RECT 207.690 70.480 208.020 70.980 ;
        RECT 207.265 70.140 208.015 70.310 ;
        RECT 207.265 69.320 207.615 69.970 ;
        RECT 207.785 69.150 208.015 70.140 ;
        RECT 207.265 68.980 208.015 69.150 ;
        RECT 201.280 68.430 206.625 68.975 ;
        RECT 207.265 68.690 207.520 68.980 ;
        RECT 207.690 68.430 208.020 68.810 ;
        RECT 208.190 68.690 208.360 70.810 ;
        RECT 208.530 70.010 208.855 70.795 ;
        RECT 209.025 70.520 209.275 70.980 ;
        RECT 209.445 70.480 209.695 70.810 ;
        RECT 209.910 70.480 210.590 70.810 ;
        RECT 209.445 70.350 209.615 70.480 ;
        RECT 209.220 70.180 209.615 70.350 ;
        RECT 208.590 68.960 209.050 70.010 ;
        RECT 209.220 68.820 209.390 70.180 ;
        RECT 209.785 69.920 210.250 70.310 ;
        RECT 209.560 69.110 209.910 69.730 ;
        RECT 210.080 69.330 210.250 69.920 ;
        RECT 210.420 69.700 210.590 70.480 ;
        RECT 210.760 70.380 210.930 70.720 ;
        RECT 211.165 70.550 211.495 70.980 ;
        RECT 211.665 70.380 211.835 70.720 ;
        RECT 212.130 70.520 212.500 70.980 ;
        RECT 210.760 70.210 211.835 70.380 ;
        RECT 212.670 70.350 212.840 70.810 ;
        RECT 213.075 70.470 213.945 70.810 ;
        RECT 214.115 70.520 214.365 70.980 ;
        RECT 212.280 70.180 212.840 70.350 ;
        RECT 212.280 70.040 212.450 70.180 ;
        RECT 210.950 69.870 212.450 70.040 ;
        RECT 213.145 70.010 213.605 70.300 ;
        RECT 210.420 69.530 212.110 69.700 ;
        RECT 210.080 69.110 210.435 69.330 ;
        RECT 210.605 68.820 210.775 69.530 ;
        RECT 210.980 69.110 211.770 69.360 ;
        RECT 211.940 69.350 212.110 69.530 ;
        RECT 212.280 69.180 212.450 69.870 ;
        RECT 208.720 68.430 209.050 68.790 ;
        RECT 209.220 68.650 209.715 68.820 ;
        RECT 209.920 68.650 210.775 68.820 ;
        RECT 211.650 68.430 211.980 68.890 ;
        RECT 212.190 68.790 212.450 69.180 ;
        RECT 212.640 70.000 213.605 70.010 ;
        RECT 213.775 70.090 213.945 70.470 ;
        RECT 214.535 70.430 214.705 70.720 ;
        RECT 214.885 70.600 215.215 70.980 ;
        RECT 214.535 70.260 215.335 70.430 ;
        RECT 212.640 69.840 213.315 70.000 ;
        RECT 213.775 69.920 214.995 70.090 ;
        RECT 212.640 69.050 212.850 69.840 ;
        RECT 213.775 69.830 213.945 69.920 ;
        RECT 213.020 69.050 213.370 69.670 ;
        RECT 213.540 69.660 213.945 69.830 ;
        RECT 213.540 68.880 213.710 69.660 ;
        RECT 213.880 69.210 214.100 69.490 ;
        RECT 214.280 69.380 214.820 69.750 ;
        RECT 215.165 69.670 215.335 70.260 ;
        RECT 215.555 69.840 215.860 70.980 ;
        RECT 216.030 69.790 216.285 70.670 ;
        RECT 215.165 69.640 215.905 69.670 ;
        RECT 213.880 69.040 214.410 69.210 ;
        RECT 212.190 68.620 212.540 68.790 ;
        RECT 212.760 68.600 213.710 68.880 ;
        RECT 213.880 68.430 214.070 68.870 ;
        RECT 214.240 68.810 214.410 69.040 ;
        RECT 214.580 68.980 214.820 69.380 ;
        RECT 214.990 69.340 215.905 69.640 ;
        RECT 214.990 69.165 215.315 69.340 ;
        RECT 214.990 68.810 215.310 69.165 ;
        RECT 216.075 69.140 216.285 69.790 ;
        RECT 216.460 70.220 216.975 70.630 ;
        RECT 217.210 70.220 217.380 70.980 ;
        RECT 217.550 70.640 219.580 70.810 ;
        RECT 216.460 69.410 216.800 70.220 ;
        RECT 217.550 69.975 217.720 70.640 ;
        RECT 218.115 70.300 219.240 70.470 ;
        RECT 216.970 69.785 217.720 69.975 ;
        RECT 217.890 69.960 218.900 70.130 ;
        RECT 216.460 69.240 217.690 69.410 ;
        RECT 214.240 68.640 215.310 68.810 ;
        RECT 215.555 68.430 215.860 68.890 ;
        RECT 216.030 68.610 216.285 69.140 ;
        RECT 216.735 68.635 216.980 69.240 ;
        RECT 217.200 68.430 217.710 68.965 ;
        RECT 217.890 68.600 218.080 69.960 ;
        RECT 218.250 68.940 218.525 69.760 ;
        RECT 218.730 69.160 218.900 69.960 ;
        RECT 219.070 69.170 219.240 70.300 ;
        RECT 219.410 69.670 219.580 70.640 ;
        RECT 219.750 69.840 219.920 70.980 ;
        RECT 220.090 69.840 220.425 70.810 ;
        RECT 220.600 70.545 225.945 70.980 ;
        RECT 219.410 69.340 219.605 69.670 ;
        RECT 219.830 69.340 220.085 69.670 ;
        RECT 219.830 69.170 220.000 69.340 ;
        RECT 220.255 69.170 220.425 69.840 ;
        RECT 219.070 69.000 220.000 69.170 ;
        RECT 219.070 68.965 219.245 69.000 ;
        RECT 218.250 68.770 218.530 68.940 ;
        RECT 218.250 68.600 218.525 68.770 ;
        RECT 218.715 68.600 219.245 68.965 ;
        RECT 219.670 68.430 220.000 68.830 ;
        RECT 220.170 68.600 220.425 69.170 ;
        RECT 222.185 68.975 222.525 69.805 ;
        RECT 224.005 69.295 224.355 70.545 ;
        RECT 226.580 69.815 226.870 70.980 ;
        RECT 227.040 70.545 232.385 70.980 ;
        RECT 220.600 68.430 225.945 68.975 ;
        RECT 226.580 68.430 226.870 69.155 ;
        RECT 228.625 68.975 228.965 69.805 ;
        RECT 230.445 69.295 230.795 70.545 ;
        RECT 232.560 69.890 234.230 70.980 ;
        RECT 232.560 69.200 233.310 69.720 ;
        RECT 233.480 69.370 234.230 69.890 ;
        RECT 234.400 70.550 234.740 70.810 ;
        RECT 227.040 68.430 232.385 68.975 ;
        RECT 232.560 68.430 234.230 69.200 ;
        RECT 234.400 69.150 234.660 70.550 ;
        RECT 234.910 70.180 235.240 70.980 ;
        RECT 235.705 70.010 235.955 70.810 ;
        RECT 236.140 70.260 236.470 70.980 ;
        RECT 236.690 70.010 236.940 70.810 ;
        RECT 237.110 70.600 237.445 70.980 ;
        RECT 234.850 69.840 237.040 70.010 ;
        RECT 234.850 69.670 235.165 69.840 ;
        RECT 234.835 69.420 235.165 69.670 ;
        RECT 234.400 68.640 234.740 69.150 ;
        RECT 234.910 68.430 235.180 69.230 ;
        RECT 235.360 68.700 235.640 69.670 ;
        RECT 235.820 68.700 236.120 69.670 ;
        RECT 236.300 68.705 236.650 69.670 ;
        RECT 236.870 68.930 237.040 69.840 ;
        RECT 237.210 69.110 237.450 70.420 ;
        RECT 237.710 70.235 237.980 70.980 ;
        RECT 238.610 70.975 244.885 70.980 ;
        RECT 238.150 70.065 238.440 70.805 ;
        RECT 238.610 70.250 238.865 70.975 ;
        RECT 239.050 70.080 239.310 70.805 ;
        RECT 239.480 70.250 239.725 70.975 ;
        RECT 239.910 70.080 240.170 70.805 ;
        RECT 240.340 70.250 240.585 70.975 ;
        RECT 240.770 70.080 241.030 70.805 ;
        RECT 241.200 70.250 241.445 70.975 ;
        RECT 241.615 70.080 241.875 70.805 ;
        RECT 242.045 70.250 242.305 70.975 ;
        RECT 242.475 70.080 242.735 70.805 ;
        RECT 242.905 70.250 243.165 70.975 ;
        RECT 243.335 70.080 243.595 70.805 ;
        RECT 243.765 70.250 244.025 70.975 ;
        RECT 244.195 70.080 244.455 70.805 ;
        RECT 244.625 70.180 244.885 70.975 ;
        RECT 239.050 70.065 244.455 70.080 ;
        RECT 237.710 69.840 244.455 70.065 ;
        RECT 237.710 69.250 238.875 69.840 ;
        RECT 245.055 69.670 245.305 70.805 ;
        RECT 245.485 70.170 245.745 70.980 ;
        RECT 245.920 69.670 246.165 70.810 ;
        RECT 246.345 70.170 246.640 70.980 ;
        RECT 246.910 69.970 247.080 70.810 ;
        RECT 247.250 70.640 248.420 70.810 ;
        RECT 247.250 70.140 247.580 70.640 ;
        RECT 248.090 70.600 248.420 70.640 ;
        RECT 248.610 70.560 248.965 70.980 ;
        RECT 247.750 70.380 247.980 70.470 ;
        RECT 249.135 70.380 249.385 70.810 ;
        RECT 247.750 70.140 249.385 70.380 ;
        RECT 249.555 70.220 249.885 70.980 ;
        RECT 250.055 70.140 250.310 70.810 ;
        RECT 246.910 69.800 249.970 69.970 ;
        RECT 239.045 69.420 246.165 69.670 ;
        RECT 237.710 69.080 244.455 69.250 ;
        RECT 236.870 68.600 237.365 68.930 ;
        RECT 237.710 68.430 238.010 68.910 ;
        RECT 238.180 68.625 238.440 69.080 ;
        RECT 238.610 68.430 238.870 68.910 ;
        RECT 239.050 68.625 239.310 69.080 ;
        RECT 239.480 68.430 239.730 68.910 ;
        RECT 239.910 68.625 240.170 69.080 ;
        RECT 240.340 68.430 240.590 68.910 ;
        RECT 240.770 68.625 241.030 69.080 ;
        RECT 241.200 68.430 241.445 68.910 ;
        RECT 241.615 68.625 241.890 69.080 ;
        RECT 242.060 68.430 242.305 68.910 ;
        RECT 242.475 68.625 242.735 69.080 ;
        RECT 242.905 68.430 243.165 68.910 ;
        RECT 243.335 68.625 243.595 69.080 ;
        RECT 243.765 68.430 244.025 68.910 ;
        RECT 244.195 68.625 244.455 69.080 ;
        RECT 244.625 68.430 244.885 68.990 ;
        RECT 245.055 68.610 245.305 69.420 ;
        RECT 245.485 68.430 245.745 68.955 ;
        RECT 245.915 68.610 246.165 69.420 ;
        RECT 246.335 69.110 246.650 69.670 ;
        RECT 246.825 69.420 247.175 69.630 ;
        RECT 247.345 69.420 247.790 69.620 ;
        RECT 247.960 69.420 248.435 69.620 ;
        RECT 246.910 69.080 247.975 69.250 ;
        RECT 246.345 68.430 246.650 68.940 ;
        RECT 246.910 68.600 247.080 69.080 ;
        RECT 247.250 68.430 247.580 68.910 ;
        RECT 247.805 68.850 247.975 69.080 ;
        RECT 248.155 69.020 248.435 69.420 ;
        RECT 248.705 69.420 249.035 69.620 ;
        RECT 249.205 69.420 249.570 69.620 ;
        RECT 248.705 69.020 248.990 69.420 ;
        RECT 249.800 69.250 249.970 69.800 ;
        RECT 249.170 69.080 249.970 69.250 ;
        RECT 249.170 68.850 249.340 69.080 ;
        RECT 250.140 69.010 250.310 70.140 ;
        RECT 250.500 69.890 252.170 70.980 ;
        RECT 250.125 68.940 250.310 69.010 ;
        RECT 250.100 68.930 250.310 68.940 ;
        RECT 247.805 68.600 249.340 68.850 ;
        RECT 249.510 68.430 249.840 68.910 ;
        RECT 250.055 68.600 250.310 68.930 ;
        RECT 250.500 69.200 251.250 69.720 ;
        RECT 251.420 69.370 252.170 69.890 ;
        RECT 252.340 69.815 252.630 70.980 ;
        RECT 252.800 69.890 256.310 70.980 ;
        RECT 252.800 69.200 254.450 69.720 ;
        RECT 254.620 69.370 256.310 69.890 ;
        RECT 257.490 69.970 257.660 70.810 ;
        RECT 257.830 70.640 259.000 70.810 ;
        RECT 257.830 70.140 258.160 70.640 ;
        RECT 258.670 70.600 259.000 70.640 ;
        RECT 259.190 70.560 259.545 70.980 ;
        RECT 258.330 70.380 258.560 70.470 ;
        RECT 259.715 70.380 259.965 70.810 ;
        RECT 258.330 70.140 259.965 70.380 ;
        RECT 260.135 70.220 260.465 70.980 ;
        RECT 260.635 70.140 260.890 70.810 ;
        RECT 257.490 69.800 260.550 69.970 ;
        RECT 257.405 69.420 257.755 69.630 ;
        RECT 257.925 69.420 258.370 69.620 ;
        RECT 258.540 69.420 259.015 69.620 ;
        RECT 250.500 68.430 252.170 69.200 ;
        RECT 252.340 68.430 252.630 69.155 ;
        RECT 252.800 68.430 256.310 69.200 ;
        RECT 257.490 69.080 258.555 69.250 ;
        RECT 257.490 68.600 257.660 69.080 ;
        RECT 257.830 68.430 258.160 68.910 ;
        RECT 258.385 68.850 258.555 69.080 ;
        RECT 258.735 69.020 259.015 69.420 ;
        RECT 259.285 69.420 259.615 69.620 ;
        RECT 259.785 69.420 260.150 69.620 ;
        RECT 259.285 69.020 259.570 69.420 ;
        RECT 260.380 69.250 260.550 69.800 ;
        RECT 259.750 69.080 260.550 69.250 ;
        RECT 259.750 68.850 259.920 69.080 ;
        RECT 260.720 69.010 260.890 70.140 ;
        RECT 261.085 70.590 261.420 70.810 ;
        RECT 262.425 70.600 262.780 70.980 ;
        RECT 261.085 69.970 261.340 70.590 ;
        RECT 261.590 70.430 261.820 70.470 ;
        RECT 262.950 70.430 263.200 70.810 ;
        RECT 261.590 70.230 263.200 70.430 ;
        RECT 261.590 70.140 261.775 70.230 ;
        RECT 262.365 70.220 263.200 70.230 ;
        RECT 263.450 70.200 263.700 70.980 ;
        RECT 263.870 70.130 264.130 70.810 ;
        RECT 264.300 70.470 265.960 70.760 ;
        RECT 261.930 70.030 262.260 70.060 ;
        RECT 261.930 69.970 263.730 70.030 ;
        RECT 261.085 69.860 263.790 69.970 ;
        RECT 261.085 69.800 262.260 69.860 ;
        RECT 263.590 69.825 263.790 69.860 ;
        RECT 261.080 69.420 261.570 69.620 ;
        RECT 261.760 69.420 262.235 69.630 ;
        RECT 260.705 68.930 260.890 69.010 ;
        RECT 258.385 68.600 259.920 68.850 ;
        RECT 260.090 68.430 260.420 68.910 ;
        RECT 260.635 68.600 260.890 68.930 ;
        RECT 261.085 68.430 261.540 69.195 ;
        RECT 262.015 69.020 262.235 69.420 ;
        RECT 262.480 69.420 262.810 69.630 ;
        RECT 262.480 69.020 262.690 69.420 ;
        RECT 262.980 69.385 263.390 69.690 ;
        RECT 263.620 69.250 263.790 69.825 ;
        RECT 263.520 69.130 263.790 69.250 ;
        RECT 262.945 69.085 263.790 69.130 ;
        RECT 262.945 68.960 263.700 69.085 ;
        RECT 262.945 68.810 263.115 68.960 ;
        RECT 263.960 68.930 264.130 70.130 ;
        RECT 264.300 70.130 265.895 70.300 ;
        RECT 266.130 70.180 266.410 70.980 ;
        RECT 264.300 69.840 264.625 70.130 ;
        RECT 265.725 70.010 265.895 70.130 ;
        RECT 264.820 69.790 265.535 69.960 ;
        RECT 265.725 69.840 266.450 70.010 ;
        RECT 266.620 69.840 266.895 70.810 ;
        RECT 264.300 69.100 264.655 69.670 ;
        RECT 264.825 69.340 265.535 69.790 ;
        RECT 266.280 69.670 266.450 69.840 ;
        RECT 265.705 69.340 266.110 69.670 ;
        RECT 266.280 69.340 266.555 69.670 ;
        RECT 266.280 69.170 266.450 69.340 ;
        RECT 264.840 69.000 266.450 69.170 ;
        RECT 266.725 69.105 266.895 69.840 ;
        RECT 267.065 69.800 267.235 70.980 ;
        RECT 267.520 70.470 268.710 70.760 ;
        RECT 267.540 70.130 268.710 70.300 ;
        RECT 268.880 70.180 269.160 70.980 ;
        RECT 267.540 69.840 267.865 70.130 ;
        RECT 268.540 70.010 268.710 70.130 ;
        RECT 268.035 69.670 268.230 69.960 ;
        RECT 268.540 69.840 269.200 70.010 ;
        RECT 269.370 69.840 269.645 70.810 ;
        RECT 269.820 69.890 271.030 70.980 ;
        RECT 271.880 70.620 272.210 70.980 ;
        RECT 272.735 70.620 273.070 70.980 ;
        RECT 273.640 70.620 273.970 70.980 ;
        RECT 274.535 70.620 274.985 70.980 ;
        RECT 269.030 69.670 269.200 69.840 ;
        RECT 261.815 68.600 263.115 68.810 ;
        RECT 263.370 68.430 263.700 68.790 ;
        RECT 263.870 68.600 264.130 68.930 ;
        RECT 264.305 68.430 264.640 68.930 ;
        RECT 264.840 68.650 265.010 69.000 ;
        RECT 265.210 68.430 265.540 68.830 ;
        RECT 265.710 68.650 265.880 69.000 ;
        RECT 266.050 68.430 266.430 68.830 ;
        RECT 266.620 68.760 266.895 69.105 ;
        RECT 267.065 68.430 267.235 69.345 ;
        RECT 267.520 69.340 267.865 69.670 ;
        RECT 268.035 69.340 268.860 69.670 ;
        RECT 269.030 69.340 269.305 69.670 ;
        RECT 269.030 69.170 269.200 69.340 ;
        RECT 267.535 69.000 269.200 69.170 ;
        RECT 269.475 69.105 269.645 69.840 ;
        RECT 267.535 68.650 267.790 69.000 ;
        RECT 267.960 68.430 268.290 68.830 ;
        RECT 268.460 68.650 268.630 69.000 ;
        RECT 268.800 68.430 269.180 68.830 ;
        RECT 269.370 68.760 269.645 69.105 ;
        RECT 269.820 69.180 270.340 69.720 ;
        RECT 270.510 69.350 271.030 69.890 ;
        RECT 271.270 70.220 275.035 70.450 ;
        RECT 269.820 68.430 271.030 69.180 ;
        RECT 271.270 68.770 271.550 70.220 ;
        RECT 271.720 68.960 272.000 70.050 ;
        RECT 272.180 69.880 273.490 70.050 ;
        RECT 272.180 69.190 272.445 69.880 ;
        RECT 273.660 69.870 274.435 70.040 ;
        RECT 273.660 69.700 273.830 69.870 ;
        RECT 272.615 69.365 273.830 69.700 ;
        RECT 272.180 68.960 273.430 69.190 ;
        RECT 273.600 69.150 273.830 69.365 ;
        RECT 274.000 69.340 274.190 69.685 ;
        RECT 273.600 68.960 274.295 69.150 ;
        RECT 274.480 69.070 274.695 69.685 ;
        RECT 274.865 69.670 275.035 70.220 ;
        RECT 275.205 69.840 275.565 70.510 ;
        RECT 275.800 69.890 277.470 70.980 ;
        RECT 274.865 69.340 275.175 69.670 ;
        RECT 275.345 69.150 275.565 69.840 ;
        RECT 271.880 68.430 272.210 68.790 ;
        RECT 272.380 68.600 272.570 68.960 ;
        RECT 273.240 68.860 273.430 68.960 ;
        RECT 274.115 68.890 274.295 68.960 ;
        RECT 275.080 68.890 275.565 69.150 ;
        RECT 272.740 68.430 273.070 68.790 ;
        RECT 273.605 68.430 273.935 68.790 ;
        RECT 274.115 68.700 275.565 68.890 ;
        RECT 275.080 68.600 275.565 68.700 ;
        RECT 275.800 69.200 276.550 69.720 ;
        RECT 276.720 69.370 277.470 69.890 ;
        RECT 278.100 69.815 278.390 70.980 ;
        RECT 278.565 70.310 278.820 70.810 ;
        RECT 278.990 70.480 279.320 70.980 ;
        RECT 278.565 70.140 279.315 70.310 ;
        RECT 278.565 69.320 278.915 69.970 ;
        RECT 275.800 68.430 277.470 69.200 ;
        RECT 278.100 68.430 278.390 69.155 ;
        RECT 279.085 69.150 279.315 70.140 ;
        RECT 278.565 68.980 279.315 69.150 ;
        RECT 278.565 68.690 278.820 68.980 ;
        RECT 278.990 68.430 279.320 68.810 ;
        RECT 279.490 68.690 279.660 70.810 ;
        RECT 279.830 70.010 280.155 70.795 ;
        RECT 280.325 70.520 280.575 70.980 ;
        RECT 280.745 70.480 280.995 70.810 ;
        RECT 281.210 70.480 281.890 70.810 ;
        RECT 280.745 70.350 280.915 70.480 ;
        RECT 280.520 70.180 280.915 70.350 ;
        RECT 279.890 68.960 280.350 70.010 ;
        RECT 280.520 68.820 280.690 70.180 ;
        RECT 281.085 69.920 281.550 70.310 ;
        RECT 280.860 69.110 281.210 69.730 ;
        RECT 281.380 69.330 281.550 69.920 ;
        RECT 281.720 69.700 281.890 70.480 ;
        RECT 282.060 70.380 282.230 70.720 ;
        RECT 282.465 70.550 282.795 70.980 ;
        RECT 282.965 70.380 283.135 70.720 ;
        RECT 283.430 70.520 283.800 70.980 ;
        RECT 282.060 70.210 283.135 70.380 ;
        RECT 283.970 70.350 284.140 70.810 ;
        RECT 284.375 70.470 285.245 70.810 ;
        RECT 285.415 70.520 285.665 70.980 ;
        RECT 283.580 70.180 284.140 70.350 ;
        RECT 283.580 70.040 283.750 70.180 ;
        RECT 282.250 69.870 283.750 70.040 ;
        RECT 284.445 70.010 284.905 70.300 ;
        RECT 281.720 69.530 283.410 69.700 ;
        RECT 281.380 69.110 281.735 69.330 ;
        RECT 281.905 68.820 282.075 69.530 ;
        RECT 282.280 69.110 283.070 69.360 ;
        RECT 283.240 69.350 283.410 69.530 ;
        RECT 283.580 69.180 283.750 69.870 ;
        RECT 280.020 68.430 280.350 68.790 ;
        RECT 280.520 68.650 281.015 68.820 ;
        RECT 281.220 68.650 282.075 68.820 ;
        RECT 282.950 68.430 283.280 68.890 ;
        RECT 283.490 68.790 283.750 69.180 ;
        RECT 283.940 70.000 284.905 70.010 ;
        RECT 285.075 70.090 285.245 70.470 ;
        RECT 285.835 70.430 286.005 70.720 ;
        RECT 286.185 70.600 286.515 70.980 ;
        RECT 285.835 70.260 286.635 70.430 ;
        RECT 283.940 69.840 284.615 70.000 ;
        RECT 285.075 69.920 286.295 70.090 ;
        RECT 283.940 69.050 284.150 69.840 ;
        RECT 285.075 69.830 285.245 69.920 ;
        RECT 284.320 69.050 284.670 69.670 ;
        RECT 284.840 69.660 285.245 69.830 ;
        RECT 284.840 68.880 285.010 69.660 ;
        RECT 285.180 69.210 285.400 69.490 ;
        RECT 285.580 69.380 286.120 69.750 ;
        RECT 286.465 69.670 286.635 70.260 ;
        RECT 286.855 69.840 287.160 70.980 ;
        RECT 287.330 69.790 287.585 70.670 ;
        RECT 286.465 69.640 287.205 69.670 ;
        RECT 285.180 69.040 285.710 69.210 ;
        RECT 283.490 68.620 283.840 68.790 ;
        RECT 284.060 68.600 285.010 68.880 ;
        RECT 285.180 68.430 285.370 68.870 ;
        RECT 285.540 68.810 285.710 69.040 ;
        RECT 285.880 68.980 286.120 69.380 ;
        RECT 286.290 69.340 287.205 69.640 ;
        RECT 286.290 69.165 286.615 69.340 ;
        RECT 286.290 68.810 286.610 69.165 ;
        RECT 287.375 69.140 287.585 69.790 ;
        RECT 285.540 68.640 286.610 68.810 ;
        RECT 286.855 68.430 287.160 68.890 ;
        RECT 287.330 68.610 287.585 69.140 ;
        RECT 288.225 69.840 288.560 70.810 ;
        RECT 288.730 69.840 288.900 70.980 ;
        RECT 289.070 70.640 291.100 70.810 ;
        RECT 288.225 69.170 288.395 69.840 ;
        RECT 289.070 69.670 289.240 70.640 ;
        RECT 288.565 69.340 288.820 69.670 ;
        RECT 289.045 69.340 289.240 69.670 ;
        RECT 289.410 70.300 290.535 70.470 ;
        RECT 288.650 69.170 288.820 69.340 ;
        RECT 289.410 69.170 289.580 70.300 ;
        RECT 288.225 68.600 288.480 69.170 ;
        RECT 288.650 69.000 289.580 69.170 ;
        RECT 289.750 69.960 290.760 70.130 ;
        RECT 289.750 69.160 289.920 69.960 ;
        RECT 289.405 68.965 289.580 69.000 ;
        RECT 288.650 68.430 288.980 68.830 ;
        RECT 289.405 68.600 289.935 68.965 ;
        RECT 290.125 68.940 290.400 69.760 ;
        RECT 290.120 68.770 290.400 68.940 ;
        RECT 290.125 68.600 290.400 68.770 ;
        RECT 290.570 68.600 290.760 69.960 ;
        RECT 290.930 69.975 291.100 70.640 ;
        RECT 291.270 70.220 291.440 70.980 ;
        RECT 291.675 70.220 292.190 70.630 ;
        RECT 290.930 69.785 291.680 69.975 ;
        RECT 291.850 69.410 292.190 70.220 ;
        RECT 292.360 69.890 294.030 70.980 ;
        RECT 294.665 70.310 294.920 70.810 ;
        RECT 295.090 70.480 295.420 70.980 ;
        RECT 294.665 70.140 295.415 70.310 ;
        RECT 290.960 69.240 292.190 69.410 ;
        RECT 290.940 68.430 291.450 68.965 ;
        RECT 291.670 68.635 291.915 69.240 ;
        RECT 292.360 69.200 293.110 69.720 ;
        RECT 293.280 69.370 294.030 69.890 ;
        RECT 294.665 69.320 295.015 69.970 ;
        RECT 292.360 68.430 294.030 69.200 ;
        RECT 295.185 69.150 295.415 70.140 ;
        RECT 294.665 68.980 295.415 69.150 ;
        RECT 294.665 68.690 294.920 68.980 ;
        RECT 295.090 68.430 295.420 68.810 ;
        RECT 295.590 68.690 295.760 70.810 ;
        RECT 295.930 70.010 296.255 70.795 ;
        RECT 296.425 70.520 296.675 70.980 ;
        RECT 296.845 70.480 297.095 70.810 ;
        RECT 297.310 70.480 297.990 70.810 ;
        RECT 296.845 70.350 297.015 70.480 ;
        RECT 296.620 70.180 297.015 70.350 ;
        RECT 295.990 68.960 296.450 70.010 ;
        RECT 296.620 68.820 296.790 70.180 ;
        RECT 297.185 69.920 297.650 70.310 ;
        RECT 296.960 69.110 297.310 69.730 ;
        RECT 297.480 69.330 297.650 69.920 ;
        RECT 297.820 69.700 297.990 70.480 ;
        RECT 298.160 70.380 298.330 70.720 ;
        RECT 298.565 70.550 298.895 70.980 ;
        RECT 299.065 70.380 299.235 70.720 ;
        RECT 299.530 70.520 299.900 70.980 ;
        RECT 298.160 70.210 299.235 70.380 ;
        RECT 300.070 70.350 300.240 70.810 ;
        RECT 300.475 70.470 301.345 70.810 ;
        RECT 301.515 70.520 301.765 70.980 ;
        RECT 299.680 70.180 300.240 70.350 ;
        RECT 299.680 70.040 299.850 70.180 ;
        RECT 298.350 69.870 299.850 70.040 ;
        RECT 300.545 70.010 301.005 70.300 ;
        RECT 297.820 69.530 299.510 69.700 ;
        RECT 297.480 69.110 297.835 69.330 ;
        RECT 298.005 68.820 298.175 69.530 ;
        RECT 298.380 69.110 299.170 69.360 ;
        RECT 299.340 69.350 299.510 69.530 ;
        RECT 299.680 69.180 299.850 69.870 ;
        RECT 296.120 68.430 296.450 68.790 ;
        RECT 296.620 68.650 297.115 68.820 ;
        RECT 297.320 68.650 298.175 68.820 ;
        RECT 299.050 68.430 299.380 68.890 ;
        RECT 299.590 68.790 299.850 69.180 ;
        RECT 300.040 70.000 301.005 70.010 ;
        RECT 301.175 70.090 301.345 70.470 ;
        RECT 301.935 70.430 302.105 70.720 ;
        RECT 302.285 70.600 302.615 70.980 ;
        RECT 301.935 70.260 302.735 70.430 ;
        RECT 300.040 69.840 300.715 70.000 ;
        RECT 301.175 69.920 302.395 70.090 ;
        RECT 300.040 69.050 300.250 69.840 ;
        RECT 301.175 69.830 301.345 69.920 ;
        RECT 300.420 69.050 300.770 69.670 ;
        RECT 300.940 69.660 301.345 69.830 ;
        RECT 300.940 68.880 301.110 69.660 ;
        RECT 301.280 69.210 301.500 69.490 ;
        RECT 301.680 69.380 302.220 69.750 ;
        RECT 302.565 69.670 302.735 70.260 ;
        RECT 302.955 69.840 303.260 70.980 ;
        RECT 303.430 69.790 303.685 70.670 ;
        RECT 303.860 69.815 304.150 70.980 ;
        RECT 304.325 69.840 304.660 70.810 ;
        RECT 304.830 69.840 305.000 70.980 ;
        RECT 305.170 70.640 307.200 70.810 ;
        RECT 302.565 69.640 303.305 69.670 ;
        RECT 301.280 69.040 301.810 69.210 ;
        RECT 299.590 68.620 299.940 68.790 ;
        RECT 300.160 68.600 301.110 68.880 ;
        RECT 301.280 68.430 301.470 68.870 ;
        RECT 301.640 68.810 301.810 69.040 ;
        RECT 301.980 68.980 302.220 69.380 ;
        RECT 302.390 69.340 303.305 69.640 ;
        RECT 302.390 69.165 302.715 69.340 ;
        RECT 302.390 68.810 302.710 69.165 ;
        RECT 303.475 69.140 303.685 69.790 ;
        RECT 304.325 69.170 304.495 69.840 ;
        RECT 305.170 69.670 305.340 70.640 ;
        RECT 304.665 69.340 304.920 69.670 ;
        RECT 305.145 69.340 305.340 69.670 ;
        RECT 305.510 70.300 306.635 70.470 ;
        RECT 304.750 69.170 304.920 69.340 ;
        RECT 305.510 69.170 305.680 70.300 ;
        RECT 301.640 68.640 302.710 68.810 ;
        RECT 302.955 68.430 303.260 68.890 ;
        RECT 303.430 68.610 303.685 69.140 ;
        RECT 303.860 68.430 304.150 69.155 ;
        RECT 304.325 68.600 304.580 69.170 ;
        RECT 304.750 69.000 305.680 69.170 ;
        RECT 305.850 69.960 306.860 70.130 ;
        RECT 305.850 69.160 306.020 69.960 ;
        RECT 306.225 69.620 306.500 69.760 ;
        RECT 306.220 69.450 306.500 69.620 ;
        RECT 305.505 68.965 305.680 69.000 ;
        RECT 304.750 68.430 305.080 68.830 ;
        RECT 305.505 68.600 306.035 68.965 ;
        RECT 306.225 68.600 306.500 69.450 ;
        RECT 306.670 68.600 306.860 69.960 ;
        RECT 307.030 69.975 307.200 70.640 ;
        RECT 307.370 70.220 307.540 70.980 ;
        RECT 307.775 70.220 308.290 70.630 ;
        RECT 307.030 69.785 307.780 69.975 ;
        RECT 307.950 69.410 308.290 70.220 ;
        RECT 307.060 69.240 308.290 69.410 ;
        RECT 308.460 69.905 308.730 70.810 ;
        RECT 308.900 70.220 309.230 70.980 ;
        RECT 309.410 70.050 309.580 70.810 ;
        RECT 307.040 68.430 307.550 68.965 ;
        RECT 307.770 68.635 308.015 69.240 ;
        RECT 308.460 69.105 308.630 69.905 ;
        RECT 308.915 69.880 309.580 70.050 ;
        RECT 309.840 69.890 311.050 70.980 ;
        RECT 308.915 69.735 309.085 69.880 ;
        RECT 308.800 69.405 309.085 69.735 ;
        RECT 308.915 69.150 309.085 69.405 ;
        RECT 309.320 69.330 309.650 69.700 ;
        RECT 309.840 69.350 310.360 69.890 ;
        RECT 310.530 69.180 311.050 69.720 ;
        RECT 308.460 68.600 308.720 69.105 ;
        RECT 308.915 68.980 309.580 69.150 ;
        RECT 308.900 68.430 309.230 68.810 ;
        RECT 309.410 68.600 309.580 68.980 ;
        RECT 309.840 68.430 311.050 69.180 ;
        RECT 162.095 68.260 311.135 68.430 ;
        RECT 162.180 67.510 163.390 68.260 ;
        RECT 162.180 66.970 162.700 67.510 ;
        RECT 163.560 67.490 167.070 68.260 ;
        RECT 167.245 67.710 167.500 68.000 ;
        RECT 167.670 67.880 168.000 68.260 ;
        RECT 167.245 67.540 167.995 67.710 ;
        RECT 162.870 66.800 163.390 67.340 ;
        RECT 163.560 66.970 165.210 67.490 ;
        RECT 165.380 66.800 167.070 67.320 ;
        RECT 162.180 65.710 163.390 66.800 ;
        RECT 163.560 65.710 167.070 66.800 ;
        RECT 167.245 66.720 167.595 67.370 ;
        RECT 167.765 66.550 167.995 67.540 ;
        RECT 167.245 66.380 167.995 66.550 ;
        RECT 167.245 65.880 167.500 66.380 ;
        RECT 167.670 65.710 168.000 66.210 ;
        RECT 168.170 65.880 168.340 68.000 ;
        RECT 168.700 67.900 169.030 68.260 ;
        RECT 169.200 67.870 169.695 68.040 ;
        RECT 169.900 67.870 170.755 68.040 ;
        RECT 168.570 66.680 169.030 67.730 ;
        RECT 168.510 65.895 168.835 66.680 ;
        RECT 169.200 66.510 169.370 67.870 ;
        RECT 169.540 66.960 169.890 67.580 ;
        RECT 170.060 67.360 170.415 67.580 ;
        RECT 170.060 66.770 170.230 67.360 ;
        RECT 170.585 67.160 170.755 67.870 ;
        RECT 171.630 67.800 171.960 68.260 ;
        RECT 172.170 67.900 172.520 68.070 ;
        RECT 170.960 67.330 171.750 67.580 ;
        RECT 172.170 67.510 172.430 67.900 ;
        RECT 172.740 67.810 173.690 68.090 ;
        RECT 173.860 67.820 174.050 68.260 ;
        RECT 174.220 67.880 175.290 68.050 ;
        RECT 171.920 67.160 172.090 67.340 ;
        RECT 169.200 66.340 169.595 66.510 ;
        RECT 169.765 66.380 170.230 66.770 ;
        RECT 170.400 66.990 172.090 67.160 ;
        RECT 169.425 66.210 169.595 66.340 ;
        RECT 170.400 66.210 170.570 66.990 ;
        RECT 172.260 66.820 172.430 67.510 ;
        RECT 170.930 66.650 172.430 66.820 ;
        RECT 172.620 66.850 172.830 67.640 ;
        RECT 173.000 67.020 173.350 67.640 ;
        RECT 173.520 67.030 173.690 67.810 ;
        RECT 174.220 67.650 174.390 67.880 ;
        RECT 173.860 67.480 174.390 67.650 ;
        RECT 173.860 67.200 174.080 67.480 ;
        RECT 174.560 67.310 174.800 67.710 ;
        RECT 173.520 66.860 173.925 67.030 ;
        RECT 174.260 66.940 174.800 67.310 ;
        RECT 174.970 67.525 175.290 67.880 ;
        RECT 175.535 67.800 175.840 68.260 ;
        RECT 176.010 67.550 176.265 68.080 ;
        RECT 174.970 67.350 175.295 67.525 ;
        RECT 174.970 67.050 175.885 67.350 ;
        RECT 175.145 67.020 175.885 67.050 ;
        RECT 172.620 66.690 173.295 66.850 ;
        RECT 173.755 66.770 173.925 66.860 ;
        RECT 172.620 66.680 173.585 66.690 ;
        RECT 172.260 66.510 172.430 66.650 ;
        RECT 169.005 65.710 169.255 66.170 ;
        RECT 169.425 65.880 169.675 66.210 ;
        RECT 169.890 65.880 170.570 66.210 ;
        RECT 170.740 66.310 171.815 66.480 ;
        RECT 172.260 66.340 172.820 66.510 ;
        RECT 173.125 66.390 173.585 66.680 ;
        RECT 173.755 66.600 174.975 66.770 ;
        RECT 170.740 65.970 170.910 66.310 ;
        RECT 171.145 65.710 171.475 66.140 ;
        RECT 171.645 65.970 171.815 66.310 ;
        RECT 172.110 65.710 172.480 66.170 ;
        RECT 172.650 65.880 172.820 66.340 ;
        RECT 173.755 66.220 173.925 66.600 ;
        RECT 175.145 66.430 175.315 67.020 ;
        RECT 176.055 66.900 176.265 67.550 ;
        RECT 176.440 67.510 177.650 68.260 ;
        RECT 177.825 67.710 178.080 68.000 ;
        RECT 178.250 67.880 178.580 68.260 ;
        RECT 177.825 67.540 178.575 67.710 ;
        RECT 176.440 66.970 176.960 67.510 ;
        RECT 173.055 65.880 173.925 66.220 ;
        RECT 174.515 66.260 175.315 66.430 ;
        RECT 174.095 65.710 174.345 66.170 ;
        RECT 174.515 65.970 174.685 66.260 ;
        RECT 174.865 65.710 175.195 66.090 ;
        RECT 175.535 65.710 175.840 66.850 ;
        RECT 176.010 66.020 176.265 66.900 ;
        RECT 177.130 66.800 177.650 67.340 ;
        RECT 176.440 65.710 177.650 66.800 ;
        RECT 177.825 66.720 178.175 67.370 ;
        RECT 178.345 66.550 178.575 67.540 ;
        RECT 177.825 66.380 178.575 66.550 ;
        RECT 177.825 65.880 178.080 66.380 ;
        RECT 178.250 65.710 178.580 66.210 ;
        RECT 178.750 65.880 178.920 68.000 ;
        RECT 179.280 67.900 179.610 68.260 ;
        RECT 179.780 67.870 180.275 68.040 ;
        RECT 180.480 67.870 181.335 68.040 ;
        RECT 179.150 66.680 179.610 67.730 ;
        RECT 179.090 65.895 179.415 66.680 ;
        RECT 179.780 66.510 179.950 67.870 ;
        RECT 180.120 66.960 180.470 67.580 ;
        RECT 180.640 67.360 180.995 67.580 ;
        RECT 180.640 66.770 180.810 67.360 ;
        RECT 181.165 67.160 181.335 67.870 ;
        RECT 182.210 67.800 182.540 68.260 ;
        RECT 182.750 67.900 183.100 68.070 ;
        RECT 181.540 67.330 182.330 67.580 ;
        RECT 182.750 67.510 183.010 67.900 ;
        RECT 183.320 67.810 184.270 68.090 ;
        RECT 184.440 67.820 184.630 68.260 ;
        RECT 184.800 67.880 185.870 68.050 ;
        RECT 182.500 67.160 182.670 67.340 ;
        RECT 179.780 66.340 180.175 66.510 ;
        RECT 180.345 66.380 180.810 66.770 ;
        RECT 180.980 66.990 182.670 67.160 ;
        RECT 180.005 66.210 180.175 66.340 ;
        RECT 180.980 66.210 181.150 66.990 ;
        RECT 182.840 66.820 183.010 67.510 ;
        RECT 181.510 66.650 183.010 66.820 ;
        RECT 183.200 66.850 183.410 67.640 ;
        RECT 183.580 67.020 183.930 67.640 ;
        RECT 184.100 67.030 184.270 67.810 ;
        RECT 184.800 67.650 184.970 67.880 ;
        RECT 184.440 67.480 184.970 67.650 ;
        RECT 184.440 67.200 184.660 67.480 ;
        RECT 185.140 67.310 185.380 67.710 ;
        RECT 184.100 66.860 184.505 67.030 ;
        RECT 184.840 66.940 185.380 67.310 ;
        RECT 185.550 67.525 185.870 67.880 ;
        RECT 186.115 67.800 186.420 68.260 ;
        RECT 186.590 67.550 186.840 68.080 ;
        RECT 185.550 67.350 185.875 67.525 ;
        RECT 185.550 67.050 186.465 67.350 ;
        RECT 185.725 67.020 186.465 67.050 ;
        RECT 183.200 66.690 183.875 66.850 ;
        RECT 184.335 66.770 184.505 66.860 ;
        RECT 183.200 66.680 184.165 66.690 ;
        RECT 182.840 66.510 183.010 66.650 ;
        RECT 179.585 65.710 179.835 66.170 ;
        RECT 180.005 65.880 180.255 66.210 ;
        RECT 180.470 65.880 181.150 66.210 ;
        RECT 181.320 66.310 182.395 66.480 ;
        RECT 182.840 66.340 183.400 66.510 ;
        RECT 183.705 66.390 184.165 66.680 ;
        RECT 184.335 66.600 185.555 66.770 ;
        RECT 181.320 65.970 181.490 66.310 ;
        RECT 181.725 65.710 182.055 66.140 ;
        RECT 182.225 65.970 182.395 66.310 ;
        RECT 182.690 65.710 183.060 66.170 ;
        RECT 183.230 65.880 183.400 66.340 ;
        RECT 184.335 66.220 184.505 66.600 ;
        RECT 185.725 66.430 185.895 67.020 ;
        RECT 186.635 66.900 186.840 67.550 ;
        RECT 187.010 67.505 187.260 68.260 ;
        RECT 187.940 67.535 188.230 68.260 ;
        RECT 188.410 67.920 189.600 68.090 ;
        RECT 188.410 67.750 188.720 67.920 ;
        RECT 188.405 66.945 188.720 67.580 ;
        RECT 183.635 65.880 184.505 66.220 ;
        RECT 185.095 66.260 185.895 66.430 ;
        RECT 184.675 65.710 184.925 66.170 ;
        RECT 185.095 65.970 185.265 66.260 ;
        RECT 185.445 65.710 185.775 66.090 ;
        RECT 186.115 65.710 186.420 66.850 ;
        RECT 186.590 66.020 186.840 66.900 ;
        RECT 187.010 65.710 187.260 66.850 ;
        RECT 187.940 65.710 188.230 66.875 ;
        RECT 188.410 65.710 188.720 66.775 ;
        RECT 188.890 66.560 189.100 67.750 ;
        RECT 189.270 67.630 189.600 67.920 ;
        RECT 189.840 67.800 190.010 68.260 ;
        RECT 190.240 67.630 190.570 68.090 ;
        RECT 190.750 67.800 190.920 68.260 ;
        RECT 191.100 67.630 191.430 68.090 ;
        RECT 189.270 67.460 191.430 67.630 ;
        RECT 191.710 67.710 191.880 68.090 ;
        RECT 192.095 67.880 192.425 68.260 ;
        RECT 191.710 67.540 192.425 67.710 ;
        RECT 189.440 66.900 189.935 67.270 ;
        RECT 190.115 67.070 190.915 67.270 ;
        RECT 191.085 66.900 191.415 67.290 ;
        RECT 191.620 66.990 191.975 67.360 ;
        RECT 192.255 67.350 192.425 67.540 ;
        RECT 192.595 67.515 192.850 68.090 ;
        RECT 192.255 67.020 192.510 67.350 ;
        RECT 189.380 66.730 191.415 66.900 ;
        RECT 192.255 66.810 192.425 67.020 ;
        RECT 191.710 66.640 192.425 66.810 ;
        RECT 192.680 66.785 192.850 67.515 ;
        RECT 193.025 67.420 193.285 68.260 ;
        RECT 193.460 67.490 196.050 68.260 ;
        RECT 193.460 66.970 194.670 67.490 ;
        RECT 196.885 67.480 197.385 68.090 ;
        RECT 188.890 66.380 190.540 66.560 ;
        RECT 188.890 65.880 189.125 66.380 ;
        RECT 190.240 66.220 190.540 66.380 ;
        RECT 189.295 65.710 189.625 66.170 ;
        RECT 189.820 66.050 190.010 66.210 ;
        RECT 190.710 66.050 190.930 66.560 ;
        RECT 189.820 65.880 190.930 66.050 ;
        RECT 191.100 65.710 191.430 66.560 ;
        RECT 191.710 65.880 191.880 66.640 ;
        RECT 192.095 65.710 192.425 66.470 ;
        RECT 192.595 65.880 192.850 66.785 ;
        RECT 193.025 65.710 193.285 66.860 ;
        RECT 194.840 66.800 196.050 67.320 ;
        RECT 196.680 67.020 197.030 67.270 ;
        RECT 197.215 66.850 197.385 67.480 ;
        RECT 198.015 67.610 198.345 68.090 ;
        RECT 198.515 67.800 198.740 68.260 ;
        RECT 198.910 67.610 199.240 68.090 ;
        RECT 198.015 67.440 199.240 67.610 ;
        RECT 199.430 67.460 199.680 68.260 ;
        RECT 199.850 67.460 200.190 68.090 ;
        RECT 200.450 67.710 200.620 68.090 ;
        RECT 200.835 67.880 201.165 68.260 ;
        RECT 200.450 67.540 201.165 67.710 ;
        RECT 197.555 67.070 197.885 67.270 ;
        RECT 198.055 67.070 198.385 67.270 ;
        RECT 198.555 67.070 198.975 67.270 ;
        RECT 199.150 67.100 199.845 67.270 ;
        RECT 199.150 66.850 199.320 67.100 ;
        RECT 200.015 66.850 200.190 67.460 ;
        RECT 200.360 66.990 200.715 67.360 ;
        RECT 200.995 67.350 201.165 67.540 ;
        RECT 201.335 67.515 201.590 68.090 ;
        RECT 200.995 67.020 201.250 67.350 ;
        RECT 193.460 65.710 196.050 66.800 ;
        RECT 196.885 66.680 199.320 66.850 ;
        RECT 196.885 65.880 197.215 66.680 ;
        RECT 197.385 65.710 197.715 66.510 ;
        RECT 198.015 65.880 198.345 66.680 ;
        RECT 198.990 65.710 199.240 66.510 ;
        RECT 199.510 65.710 199.680 66.850 ;
        RECT 199.850 65.880 200.190 66.850 ;
        RECT 200.995 66.810 201.165 67.020 ;
        RECT 200.450 66.640 201.165 66.810 ;
        RECT 201.420 66.785 201.590 67.515 ;
        RECT 201.765 67.420 202.025 68.260 ;
        RECT 202.200 67.715 207.545 68.260 ;
        RECT 203.785 66.885 204.125 67.715 ;
        RECT 207.720 67.630 208.060 68.090 ;
        RECT 208.230 67.800 208.400 68.260 ;
        RECT 209.030 67.825 209.390 68.090 ;
        RECT 209.035 67.820 209.390 67.825 ;
        RECT 209.040 67.810 209.390 67.820 ;
        RECT 209.045 67.805 209.390 67.810 ;
        RECT 209.050 67.795 209.390 67.805 ;
        RECT 209.630 67.800 209.800 68.260 ;
        RECT 209.055 67.790 209.390 67.795 ;
        RECT 209.065 67.780 209.390 67.790 ;
        RECT 209.075 67.770 209.390 67.780 ;
        RECT 208.570 67.630 208.900 67.710 ;
        RECT 207.720 67.440 208.900 67.630 ;
        RECT 209.090 67.630 209.390 67.770 ;
        RECT 209.090 67.440 209.800 67.630 ;
        RECT 200.450 65.880 200.620 66.640 ;
        RECT 200.835 65.710 201.165 66.470 ;
        RECT 201.335 65.880 201.590 66.785 ;
        RECT 201.765 65.710 202.025 66.860 ;
        RECT 205.605 66.145 205.955 67.395 ;
        RECT 207.720 67.070 208.050 67.270 ;
        RECT 208.360 67.250 208.690 67.270 ;
        RECT 208.240 67.070 208.690 67.250 ;
        RECT 207.720 66.730 207.950 67.070 ;
        RECT 202.200 65.710 207.545 66.145 ;
        RECT 207.730 65.710 208.060 66.430 ;
        RECT 208.240 65.955 208.455 67.070 ;
        RECT 208.860 67.040 209.330 67.270 ;
        RECT 209.515 66.870 209.800 67.440 ;
        RECT 209.970 67.315 210.310 68.090 ;
        RECT 210.810 67.860 211.140 68.260 ;
        RECT 211.310 67.690 211.640 68.030 ;
        RECT 212.690 67.860 213.020 68.260 ;
        RECT 208.650 66.655 209.800 66.870 ;
        RECT 208.650 65.880 208.980 66.655 ;
        RECT 209.150 65.710 209.860 66.485 ;
        RECT 210.030 65.880 210.310 67.315 ;
        RECT 210.655 67.520 213.020 67.690 ;
        RECT 213.190 67.535 213.520 68.045 ;
        RECT 213.700 67.535 213.990 68.260 ;
        RECT 210.655 66.520 210.825 67.520 ;
        RECT 212.850 67.350 213.020 67.520 ;
        RECT 210.995 66.690 211.240 67.350 ;
        RECT 211.455 66.690 211.720 67.350 ;
        RECT 211.915 66.690 212.200 67.350 ;
        RECT 212.375 67.020 212.680 67.350 ;
        RECT 212.850 67.020 213.160 67.350 ;
        RECT 212.375 66.690 212.590 67.020 ;
        RECT 210.655 66.350 211.110 66.520 ;
        RECT 210.780 65.920 211.110 66.350 ;
        RECT 211.290 66.350 212.580 66.520 ;
        RECT 211.290 65.930 211.540 66.350 ;
        RECT 211.770 65.710 212.100 66.180 ;
        RECT 212.330 65.930 212.580 66.350 ;
        RECT 212.770 65.710 213.020 66.850 ;
        RECT 213.330 66.770 213.520 67.535 ;
        RECT 214.365 67.480 214.865 68.090 ;
        RECT 214.160 67.020 214.510 67.270 ;
        RECT 213.190 65.920 213.520 66.770 ;
        RECT 213.700 65.710 213.990 66.875 ;
        RECT 214.695 66.850 214.865 67.480 ;
        RECT 215.495 67.610 215.825 68.090 ;
        RECT 215.995 67.800 216.220 68.260 ;
        RECT 216.390 67.610 216.720 68.090 ;
        RECT 215.495 67.440 216.720 67.610 ;
        RECT 216.910 67.460 217.160 68.260 ;
        RECT 217.330 67.460 217.670 68.090 ;
        RECT 217.845 67.495 218.300 68.260 ;
        RECT 218.575 67.880 219.875 68.090 ;
        RECT 220.130 67.900 220.460 68.260 ;
        RECT 219.705 67.730 219.875 67.880 ;
        RECT 220.630 67.760 220.890 68.090 ;
        RECT 215.035 67.070 215.365 67.270 ;
        RECT 215.535 67.070 215.865 67.270 ;
        RECT 216.035 67.070 216.455 67.270 ;
        RECT 216.630 67.100 217.325 67.270 ;
        RECT 216.630 66.850 216.800 67.100 ;
        RECT 217.495 66.850 217.670 67.460 ;
        RECT 218.775 67.270 218.995 67.670 ;
        RECT 217.840 67.070 218.330 67.270 ;
        RECT 218.520 67.060 218.995 67.270 ;
        RECT 219.240 67.270 219.450 67.670 ;
        RECT 219.705 67.605 220.460 67.730 ;
        RECT 219.705 67.560 220.550 67.605 ;
        RECT 220.280 67.440 220.550 67.560 ;
        RECT 219.240 67.060 219.570 67.270 ;
        RECT 219.740 67.000 220.150 67.305 ;
        RECT 214.365 66.680 216.800 66.850 ;
        RECT 214.365 65.880 214.695 66.680 ;
        RECT 214.865 65.710 215.195 66.510 ;
        RECT 215.495 65.880 215.825 66.680 ;
        RECT 216.470 65.710 216.720 66.510 ;
        RECT 216.990 65.710 217.160 66.850 ;
        RECT 217.330 65.880 217.670 66.850 ;
        RECT 217.845 66.830 219.020 66.890 ;
        RECT 220.380 66.865 220.550 67.440 ;
        RECT 220.350 66.830 220.550 66.865 ;
        RECT 217.845 66.720 220.550 66.830 ;
        RECT 217.845 66.100 218.100 66.720 ;
        RECT 218.690 66.660 220.490 66.720 ;
        RECT 218.690 66.630 219.020 66.660 ;
        RECT 220.720 66.560 220.890 67.760 ;
        RECT 221.060 67.490 224.570 68.260 ;
        RECT 224.740 67.510 225.950 68.260 ;
        RECT 226.120 67.880 227.505 68.090 ;
        RECT 226.120 67.610 226.410 67.880 ;
        RECT 226.580 67.520 227.005 67.710 ;
        RECT 227.175 67.690 227.505 67.880 ;
        RECT 227.740 67.860 228.070 68.260 ;
        RECT 228.245 67.690 228.575 68.090 ;
        RECT 228.780 67.700 228.950 68.260 ;
        RECT 227.175 67.520 228.575 67.690 ;
        RECT 229.120 67.520 229.630 68.090 ;
        RECT 221.060 66.970 222.710 67.490 ;
        RECT 222.880 66.800 224.570 67.320 ;
        RECT 224.740 66.970 225.260 67.510 ;
        RECT 225.430 66.800 225.950 67.340 ;
        RECT 226.120 67.020 226.395 67.350 ;
        RECT 218.350 66.460 218.535 66.550 ;
        RECT 219.125 66.460 219.960 66.470 ;
        RECT 218.350 66.260 219.960 66.460 ;
        RECT 218.350 66.220 218.580 66.260 ;
        RECT 217.845 65.880 218.180 66.100 ;
        RECT 219.185 65.710 219.540 66.090 ;
        RECT 219.710 65.880 219.960 66.260 ;
        RECT 220.210 65.710 220.460 66.490 ;
        RECT 220.630 65.880 220.890 66.560 ;
        RECT 221.060 65.710 224.570 66.800 ;
        RECT 224.740 65.710 225.950 66.800 ;
        RECT 226.120 65.710 226.410 66.850 ;
        RECT 226.580 66.510 226.750 67.520 ;
        RECT 226.920 66.685 227.275 67.350 ;
        RECT 227.460 66.685 227.735 67.350 ;
        RECT 227.905 67.020 228.250 67.350 ;
        RECT 228.540 67.270 228.710 67.350 ;
        RECT 229.080 67.270 229.270 67.350 ;
        RECT 228.460 67.020 228.710 67.270 ;
        RECT 228.905 67.020 229.270 67.270 ;
        RECT 226.580 66.260 227.535 66.510 ;
        RECT 227.205 66.050 227.535 66.260 ;
        RECT 227.905 66.220 228.230 67.020 ;
        RECT 228.905 66.850 229.075 67.020 ;
        RECT 229.455 66.850 229.630 67.520 ;
        RECT 229.800 67.510 231.010 68.260 ;
        RECT 231.180 67.800 231.740 68.090 ;
        RECT 231.910 67.800 232.160 68.260 ;
        RECT 229.800 66.970 230.320 67.510 ;
        RECT 228.400 66.680 229.075 66.850 ;
        RECT 228.400 66.050 228.570 66.680 ;
        RECT 227.205 65.880 228.570 66.050 ;
        RECT 228.740 65.710 229.030 66.510 ;
        RECT 229.245 65.890 229.630 66.850 ;
        RECT 230.490 66.800 231.010 67.340 ;
        RECT 229.800 65.710 231.010 66.800 ;
        RECT 231.180 66.430 231.430 67.800 ;
        RECT 232.780 67.630 233.110 67.990 ;
        RECT 233.480 67.715 238.825 68.260 ;
        RECT 231.720 67.440 233.110 67.630 ;
        RECT 231.720 67.350 231.890 67.440 ;
        RECT 231.600 67.020 231.890 67.350 ;
        RECT 232.060 67.020 232.400 67.270 ;
        RECT 232.620 67.020 233.295 67.270 ;
        RECT 231.720 66.770 231.890 67.020 ;
        RECT 231.720 66.600 232.660 66.770 ;
        RECT 233.030 66.660 233.295 67.020 ;
        RECT 235.065 66.885 235.405 67.715 ;
        RECT 239.460 67.535 239.750 68.260 ;
        RECT 239.925 67.585 240.200 67.930 ;
        RECT 240.390 67.860 240.770 68.260 ;
        RECT 240.940 67.690 241.110 68.040 ;
        RECT 241.280 67.860 241.610 68.260 ;
        RECT 241.780 67.690 242.035 68.040 ;
        RECT 231.180 65.880 231.640 66.430 ;
        RECT 231.830 65.710 232.160 66.430 ;
        RECT 232.360 66.050 232.660 66.600 ;
        RECT 232.830 65.710 233.110 66.380 ;
        RECT 236.885 66.145 237.235 67.395 ;
        RECT 233.480 65.710 238.825 66.145 ;
        RECT 239.460 65.710 239.750 66.875 ;
        RECT 239.925 66.850 240.095 67.585 ;
        RECT 240.370 67.520 242.035 67.690 ;
        RECT 240.370 67.350 240.540 67.520 ;
        RECT 240.265 67.020 240.540 67.350 ;
        RECT 240.710 67.020 241.535 67.350 ;
        RECT 241.705 67.020 242.050 67.350 ;
        RECT 240.370 66.850 240.540 67.020 ;
        RECT 239.925 65.880 240.200 66.850 ;
        RECT 240.370 66.680 241.030 66.850 ;
        RECT 241.340 66.730 241.535 67.020 ;
        RECT 240.860 66.560 241.030 66.680 ;
        RECT 241.705 66.560 242.030 66.850 ;
        RECT 240.410 65.710 240.690 66.510 ;
        RECT 240.860 66.390 242.030 66.560 ;
        RECT 240.860 65.930 242.050 66.220 ;
        RECT 242.220 65.880 242.480 68.090 ;
        RECT 242.650 67.880 242.980 68.260 ;
        RECT 243.190 67.350 243.385 67.925 ;
        RECT 243.655 67.350 243.840 67.930 ;
        RECT 242.650 66.430 242.820 67.350 ;
        RECT 243.130 67.020 243.385 67.350 ;
        RECT 243.610 67.020 243.840 67.350 ;
        RECT 244.090 67.920 245.570 68.090 ;
        RECT 244.090 67.020 244.260 67.920 ;
        RECT 244.430 67.420 244.980 67.750 ;
        RECT 245.170 67.590 245.570 67.920 ;
        RECT 245.750 67.880 246.080 68.260 ;
        RECT 246.390 67.760 246.650 68.090 ;
        RECT 243.190 66.710 243.385 67.020 ;
        RECT 243.655 66.710 243.840 67.020 ;
        RECT 244.430 66.430 244.600 67.420 ;
        RECT 245.170 67.110 245.340 67.590 ;
        RECT 245.920 67.400 246.130 67.580 ;
        RECT 245.510 67.230 246.130 67.400 ;
        RECT 242.650 66.260 244.600 66.430 ;
        RECT 244.770 66.940 245.340 67.110 ;
        RECT 246.480 67.060 246.650 67.760 ;
        RECT 246.820 67.715 252.165 68.260 ;
        RECT 252.340 67.715 257.685 68.260 ;
        RECT 244.770 66.430 244.940 66.940 ;
        RECT 245.520 66.890 246.650 67.060 ;
        RECT 245.520 66.770 245.690 66.890 ;
        RECT 245.110 66.600 245.690 66.770 ;
        RECT 244.770 66.260 245.510 66.430 ;
        RECT 245.960 66.390 246.310 66.720 ;
        RECT 242.650 65.710 242.980 66.090 ;
        RECT 243.405 65.880 243.575 66.260 ;
        RECT 243.835 65.710 244.165 66.090 ;
        RECT 244.360 65.880 244.530 66.260 ;
        RECT 244.740 65.710 245.070 66.090 ;
        RECT 245.320 65.880 245.510 66.260 ;
        RECT 246.480 66.210 246.650 66.890 ;
        RECT 248.405 66.885 248.745 67.715 ;
        RECT 245.750 65.710 246.080 66.090 ;
        RECT 246.390 65.880 246.650 66.210 ;
        RECT 250.225 66.145 250.575 67.395 ;
        RECT 253.925 66.885 254.265 67.715 ;
        RECT 257.860 67.490 261.370 68.260 ;
        RECT 262.200 67.630 262.530 67.990 ;
        RECT 263.150 67.800 263.400 68.260 ;
        RECT 263.570 67.800 264.130 68.090 ;
        RECT 255.745 66.145 256.095 67.395 ;
        RECT 257.860 66.970 259.510 67.490 ;
        RECT 262.200 67.440 263.590 67.630 ;
        RECT 263.420 67.350 263.590 67.440 ;
        RECT 259.680 66.800 261.370 67.320 ;
        RECT 246.820 65.710 252.165 66.145 ;
        RECT 252.340 65.710 257.685 66.145 ;
        RECT 257.860 65.710 261.370 66.800 ;
        RECT 262.015 67.020 262.690 67.270 ;
        RECT 262.910 67.020 263.250 67.270 ;
        RECT 263.420 67.020 263.710 67.350 ;
        RECT 262.015 66.660 262.280 67.020 ;
        RECT 263.420 66.770 263.590 67.020 ;
        RECT 262.650 66.600 263.590 66.770 ;
        RECT 262.200 65.710 262.480 66.380 ;
        RECT 262.650 66.050 262.950 66.600 ;
        RECT 263.880 66.430 264.130 67.800 ;
        RECT 265.220 67.535 265.510 68.260 ;
        RECT 265.680 67.715 271.025 68.260 ;
        RECT 267.265 66.885 267.605 67.715 ;
        RECT 272.125 67.440 272.400 68.260 ;
        RECT 272.570 67.620 272.900 68.090 ;
        RECT 273.070 67.790 273.240 68.260 ;
        RECT 273.410 67.620 273.740 68.090 ;
        RECT 273.910 67.790 274.200 68.260 ;
        RECT 274.420 67.715 279.765 68.260 ;
        RECT 272.570 67.610 273.740 67.620 ;
        RECT 272.570 67.580 274.170 67.610 ;
        RECT 272.570 67.440 274.190 67.580 ;
        RECT 273.955 67.410 274.190 67.440 ;
        RECT 263.150 65.710 263.480 66.430 ;
        RECT 263.670 65.880 264.130 66.430 ;
        RECT 265.220 65.710 265.510 66.875 ;
        RECT 269.085 66.145 269.435 67.395 ;
        RECT 272.125 67.070 272.845 67.270 ;
        RECT 273.015 67.070 273.785 67.270 ;
        RECT 273.955 66.900 274.170 67.410 ;
        RECT 272.125 66.680 273.240 66.890 ;
        RECT 265.680 65.710 271.025 66.145 ;
        RECT 272.125 65.880 272.400 66.680 ;
        RECT 272.570 65.710 272.900 66.510 ;
        RECT 273.070 66.050 273.240 66.680 ;
        RECT 273.410 66.680 274.170 66.900 ;
        RECT 276.005 66.885 276.345 67.715 ;
        RECT 279.945 67.520 280.200 68.090 ;
        RECT 280.370 67.860 280.700 68.260 ;
        RECT 281.125 67.725 281.655 68.090 ;
        RECT 281.125 67.690 281.300 67.725 ;
        RECT 280.370 67.520 281.300 67.690 ;
        RECT 273.410 66.220 273.740 66.680 ;
        RECT 273.910 66.050 274.210 66.510 ;
        RECT 277.825 66.145 278.175 67.395 ;
        RECT 279.945 66.850 280.115 67.520 ;
        RECT 280.370 67.350 280.540 67.520 ;
        RECT 280.285 67.020 280.540 67.350 ;
        RECT 280.765 67.020 280.960 67.350 ;
        RECT 273.070 65.880 274.210 66.050 ;
        RECT 274.420 65.710 279.765 66.145 ;
        RECT 279.945 65.880 280.280 66.850 ;
        RECT 280.450 65.710 280.620 66.850 ;
        RECT 280.790 66.050 280.960 67.020 ;
        RECT 281.130 66.390 281.300 67.520 ;
        RECT 281.470 66.730 281.640 67.530 ;
        RECT 281.845 67.240 282.120 68.090 ;
        RECT 281.840 67.070 282.120 67.240 ;
        RECT 281.845 66.930 282.120 67.070 ;
        RECT 282.290 66.730 282.480 68.090 ;
        RECT 282.660 67.725 283.170 68.260 ;
        RECT 283.390 67.450 283.635 68.055 ;
        RECT 284.080 67.630 284.420 68.090 ;
        RECT 284.590 67.800 284.760 68.260 ;
        RECT 285.390 67.825 285.750 68.090 ;
        RECT 285.395 67.820 285.750 67.825 ;
        RECT 285.400 67.810 285.750 67.820 ;
        RECT 285.405 67.805 285.750 67.810 ;
        RECT 285.410 67.795 285.750 67.805 ;
        RECT 285.990 67.800 286.160 68.260 ;
        RECT 285.415 67.790 285.750 67.795 ;
        RECT 285.425 67.780 285.750 67.790 ;
        RECT 285.435 67.770 285.750 67.780 ;
        RECT 284.930 67.630 285.260 67.710 ;
        RECT 282.680 67.280 283.910 67.450 ;
        RECT 284.080 67.440 285.260 67.630 ;
        RECT 285.450 67.630 285.750 67.770 ;
        RECT 285.450 67.440 286.160 67.630 ;
        RECT 281.470 66.560 282.480 66.730 ;
        RECT 282.650 66.715 283.400 66.905 ;
        RECT 281.130 66.220 282.255 66.390 ;
        RECT 282.650 66.050 282.820 66.715 ;
        RECT 283.570 66.470 283.910 67.280 ;
        RECT 284.080 67.070 284.410 67.270 ;
        RECT 284.720 67.250 285.050 67.270 ;
        RECT 284.600 67.070 285.050 67.250 ;
        RECT 284.080 66.730 284.310 67.070 ;
        RECT 280.790 65.880 282.820 66.050 ;
        RECT 282.990 65.710 283.160 66.470 ;
        RECT 283.395 66.060 283.910 66.470 ;
        RECT 284.090 65.710 284.420 66.430 ;
        RECT 284.600 65.955 284.815 67.070 ;
        RECT 285.220 67.040 285.690 67.270 ;
        RECT 285.875 66.870 286.160 67.440 ;
        RECT 286.330 67.315 286.670 68.090 ;
        RECT 285.010 66.655 286.160 66.870 ;
        RECT 285.010 65.880 285.340 66.655 ;
        RECT 285.510 65.710 286.220 66.485 ;
        RECT 286.390 65.880 286.670 67.315 ;
        RECT 286.840 67.490 290.350 68.260 ;
        RECT 290.980 67.535 291.270 68.260 ;
        RECT 291.440 67.490 294.950 68.260 ;
        RECT 295.125 67.520 295.380 68.090 ;
        RECT 295.550 67.860 295.880 68.260 ;
        RECT 296.305 67.725 296.835 68.090 ;
        RECT 296.305 67.690 296.480 67.725 ;
        RECT 295.550 67.520 296.480 67.690 ;
        RECT 297.025 67.580 297.300 68.090 ;
        RECT 286.840 66.970 288.490 67.490 ;
        RECT 288.660 66.800 290.350 67.320 ;
        RECT 291.440 66.970 293.090 67.490 ;
        RECT 286.840 65.710 290.350 66.800 ;
        RECT 290.980 65.710 291.270 66.875 ;
        RECT 293.260 66.800 294.950 67.320 ;
        RECT 291.440 65.710 294.950 66.800 ;
        RECT 295.125 66.850 295.295 67.520 ;
        RECT 295.550 67.350 295.720 67.520 ;
        RECT 295.465 67.020 295.720 67.350 ;
        RECT 295.945 67.020 296.140 67.350 ;
        RECT 295.125 65.880 295.460 66.850 ;
        RECT 295.630 65.710 295.800 66.850 ;
        RECT 295.970 66.050 296.140 67.020 ;
        RECT 296.310 66.390 296.480 67.520 ;
        RECT 296.650 66.730 296.820 67.530 ;
        RECT 297.020 67.410 297.300 67.580 ;
        RECT 297.025 66.930 297.300 67.410 ;
        RECT 297.470 66.730 297.660 68.090 ;
        RECT 297.840 67.725 298.350 68.260 ;
        RECT 298.570 67.450 298.815 68.055 ;
        RECT 299.265 67.710 299.520 68.000 ;
        RECT 299.690 67.880 300.020 68.260 ;
        RECT 299.265 67.540 300.015 67.710 ;
        RECT 297.860 67.280 299.090 67.450 ;
        RECT 296.650 66.560 297.660 66.730 ;
        RECT 297.830 66.715 298.580 66.905 ;
        RECT 296.310 66.220 297.435 66.390 ;
        RECT 297.830 66.050 298.000 66.715 ;
        RECT 298.750 66.470 299.090 67.280 ;
        RECT 299.265 66.720 299.615 67.370 ;
        RECT 299.785 66.550 300.015 67.540 ;
        RECT 295.970 65.880 298.000 66.050 ;
        RECT 298.170 65.710 298.340 66.470 ;
        RECT 298.575 66.060 299.090 66.470 ;
        RECT 299.265 66.380 300.015 66.550 ;
        RECT 299.265 65.880 299.520 66.380 ;
        RECT 299.690 65.710 300.020 66.210 ;
        RECT 300.190 65.880 300.360 68.000 ;
        RECT 300.720 67.900 301.050 68.260 ;
        RECT 301.220 67.870 301.715 68.040 ;
        RECT 301.920 67.870 302.775 68.040 ;
        RECT 300.590 66.680 301.050 67.730 ;
        RECT 300.530 65.895 300.855 66.680 ;
        RECT 301.220 66.510 301.390 67.870 ;
        RECT 301.560 66.960 301.910 67.580 ;
        RECT 302.080 67.360 302.435 67.580 ;
        RECT 302.080 66.770 302.250 67.360 ;
        RECT 302.605 67.160 302.775 67.870 ;
        RECT 303.650 67.800 303.980 68.260 ;
        RECT 304.190 67.900 304.540 68.070 ;
        RECT 302.980 67.330 303.770 67.580 ;
        RECT 304.190 67.510 304.450 67.900 ;
        RECT 304.760 67.810 305.710 68.090 ;
        RECT 305.880 67.820 306.070 68.260 ;
        RECT 306.240 67.880 307.310 68.050 ;
        RECT 303.940 67.160 304.110 67.340 ;
        RECT 301.220 66.340 301.615 66.510 ;
        RECT 301.785 66.380 302.250 66.770 ;
        RECT 302.420 66.990 304.110 67.160 ;
        RECT 301.445 66.210 301.615 66.340 ;
        RECT 302.420 66.210 302.590 66.990 ;
        RECT 304.280 66.820 304.450 67.510 ;
        RECT 302.950 66.650 304.450 66.820 ;
        RECT 304.640 66.850 304.850 67.640 ;
        RECT 305.020 67.020 305.370 67.640 ;
        RECT 305.540 67.030 305.710 67.810 ;
        RECT 306.240 67.650 306.410 67.880 ;
        RECT 305.880 67.480 306.410 67.650 ;
        RECT 305.880 67.200 306.100 67.480 ;
        RECT 306.580 67.310 306.820 67.710 ;
        RECT 305.540 66.860 305.945 67.030 ;
        RECT 306.280 66.940 306.820 67.310 ;
        RECT 306.990 67.525 307.310 67.880 ;
        RECT 307.555 67.800 307.860 68.260 ;
        RECT 308.030 67.550 308.280 68.080 ;
        RECT 306.990 67.350 307.315 67.525 ;
        RECT 306.990 67.050 307.905 67.350 ;
        RECT 307.165 67.020 307.905 67.050 ;
        RECT 304.640 66.690 305.315 66.850 ;
        RECT 305.775 66.770 305.945 66.860 ;
        RECT 304.640 66.680 305.605 66.690 ;
        RECT 304.280 66.510 304.450 66.650 ;
        RECT 301.025 65.710 301.275 66.170 ;
        RECT 301.445 65.880 301.695 66.210 ;
        RECT 301.910 65.880 302.590 66.210 ;
        RECT 302.760 66.310 303.835 66.480 ;
        RECT 304.280 66.340 304.840 66.510 ;
        RECT 305.145 66.390 305.605 66.680 ;
        RECT 305.775 66.600 306.995 66.770 ;
        RECT 302.760 65.970 302.930 66.310 ;
        RECT 303.165 65.710 303.495 66.140 ;
        RECT 303.665 65.970 303.835 66.310 ;
        RECT 304.130 65.710 304.500 66.170 ;
        RECT 304.670 65.880 304.840 66.340 ;
        RECT 305.775 66.220 305.945 66.600 ;
        RECT 307.165 66.430 307.335 67.020 ;
        RECT 308.075 66.900 308.280 67.550 ;
        RECT 308.450 67.505 308.700 68.260 ;
        RECT 309.840 67.510 311.050 68.260 ;
        RECT 305.075 65.880 305.945 66.220 ;
        RECT 306.535 66.260 307.335 66.430 ;
        RECT 306.115 65.710 306.365 66.170 ;
        RECT 306.535 65.970 306.705 66.260 ;
        RECT 306.885 65.710 307.215 66.090 ;
        RECT 307.555 65.710 307.860 66.850 ;
        RECT 308.030 66.020 308.280 66.900 ;
        RECT 308.450 65.710 308.700 66.850 ;
        RECT 309.840 66.800 310.360 67.340 ;
        RECT 310.530 66.970 311.050 67.510 ;
        RECT 309.840 65.710 311.050 66.800 ;
        RECT 162.095 65.540 311.135 65.710 ;
        RECT 162.180 64.450 163.390 65.540 ;
        RECT 163.560 64.450 165.230 65.540 ;
        RECT 162.180 63.740 162.700 64.280 ;
        RECT 162.870 63.910 163.390 64.450 ;
        RECT 163.560 63.760 164.310 64.280 ;
        RECT 164.480 63.930 165.230 64.450 ;
        RECT 165.450 64.400 165.700 65.540 ;
        RECT 165.870 64.350 166.120 65.230 ;
        RECT 166.290 64.400 166.595 65.540 ;
        RECT 166.935 65.160 167.265 65.540 ;
        RECT 167.445 64.990 167.615 65.280 ;
        RECT 167.785 65.080 168.035 65.540 ;
        RECT 166.815 64.820 167.615 64.990 ;
        RECT 168.205 65.030 169.075 65.370 ;
        RECT 162.180 62.990 163.390 63.740 ;
        RECT 163.560 62.990 165.230 63.760 ;
        RECT 165.450 62.990 165.700 63.745 ;
        RECT 165.870 63.700 166.075 64.350 ;
        RECT 166.815 64.230 166.985 64.820 ;
        RECT 168.205 64.650 168.375 65.030 ;
        RECT 169.310 64.910 169.480 65.370 ;
        RECT 169.650 65.080 170.020 65.540 ;
        RECT 170.315 64.940 170.485 65.280 ;
        RECT 170.655 65.110 170.985 65.540 ;
        RECT 171.220 64.940 171.390 65.280 ;
        RECT 167.155 64.480 168.375 64.650 ;
        RECT 168.545 64.570 169.005 64.860 ;
        RECT 169.310 64.740 169.870 64.910 ;
        RECT 170.315 64.770 171.390 64.940 ;
        RECT 171.560 65.040 172.240 65.370 ;
        RECT 172.455 65.040 172.705 65.370 ;
        RECT 172.875 65.080 173.125 65.540 ;
        RECT 169.700 64.600 169.870 64.740 ;
        RECT 168.545 64.560 169.510 64.570 ;
        RECT 168.205 64.390 168.375 64.480 ;
        RECT 168.835 64.400 169.510 64.560 ;
        RECT 166.245 64.200 166.985 64.230 ;
        RECT 166.245 63.900 167.160 64.200 ;
        RECT 166.835 63.725 167.160 63.900 ;
        RECT 165.870 63.170 166.120 63.700 ;
        RECT 166.290 62.990 166.595 63.450 ;
        RECT 166.840 63.370 167.160 63.725 ;
        RECT 167.330 63.940 167.870 64.310 ;
        RECT 168.205 64.220 168.610 64.390 ;
        RECT 167.330 63.540 167.570 63.940 ;
        RECT 168.050 63.770 168.270 64.050 ;
        RECT 167.740 63.600 168.270 63.770 ;
        RECT 167.740 63.370 167.910 63.600 ;
        RECT 168.440 63.440 168.610 64.220 ;
        RECT 168.780 63.610 169.130 64.230 ;
        RECT 169.300 63.610 169.510 64.400 ;
        RECT 169.700 64.430 171.200 64.600 ;
        RECT 169.700 63.740 169.870 64.430 ;
        RECT 171.560 64.260 171.730 65.040 ;
        RECT 172.535 64.910 172.705 65.040 ;
        RECT 170.040 64.090 171.730 64.260 ;
        RECT 171.900 64.480 172.365 64.870 ;
        RECT 172.535 64.740 172.930 64.910 ;
        RECT 170.040 63.910 170.210 64.090 ;
        RECT 166.840 63.200 167.910 63.370 ;
        RECT 168.080 62.990 168.270 63.430 ;
        RECT 168.440 63.160 169.390 63.440 ;
        RECT 169.700 63.350 169.960 63.740 ;
        RECT 170.380 63.670 171.170 63.920 ;
        RECT 169.610 63.180 169.960 63.350 ;
        RECT 170.170 62.990 170.500 63.450 ;
        RECT 171.375 63.380 171.545 64.090 ;
        RECT 171.900 63.890 172.070 64.480 ;
        RECT 171.715 63.670 172.070 63.890 ;
        RECT 172.240 63.670 172.590 64.290 ;
        RECT 172.760 63.380 172.930 64.740 ;
        RECT 173.295 64.570 173.620 65.355 ;
        RECT 173.100 63.520 173.560 64.570 ;
        RECT 171.375 63.210 172.230 63.380 ;
        RECT 172.435 63.210 172.930 63.380 ;
        RECT 173.100 62.990 173.430 63.350 ;
        RECT 173.790 63.250 173.960 65.370 ;
        RECT 174.130 65.040 174.460 65.540 ;
        RECT 174.630 64.870 174.885 65.370 ;
        RECT 174.135 64.700 174.885 64.870 ;
        RECT 174.135 63.710 174.365 64.700 ;
        RECT 174.535 63.880 174.885 64.530 ;
        RECT 175.060 64.375 175.350 65.540 ;
        RECT 175.525 64.400 175.860 65.370 ;
        RECT 176.030 64.400 176.200 65.540 ;
        RECT 176.370 65.200 178.400 65.370 ;
        RECT 175.525 63.730 175.695 64.400 ;
        RECT 176.370 64.230 176.540 65.200 ;
        RECT 175.865 63.900 176.120 64.230 ;
        RECT 176.345 63.900 176.540 64.230 ;
        RECT 176.710 64.860 177.835 65.030 ;
        RECT 175.950 63.730 176.120 63.900 ;
        RECT 176.710 63.730 176.880 64.860 ;
        RECT 174.135 63.540 174.885 63.710 ;
        RECT 174.130 62.990 174.460 63.370 ;
        RECT 174.630 63.250 174.885 63.540 ;
        RECT 175.060 62.990 175.350 63.715 ;
        RECT 175.525 63.160 175.780 63.730 ;
        RECT 175.950 63.560 176.880 63.730 ;
        RECT 177.050 64.520 178.060 64.690 ;
        RECT 177.050 63.720 177.220 64.520 ;
        RECT 177.425 64.180 177.700 64.320 ;
        RECT 177.420 64.010 177.700 64.180 ;
        RECT 176.705 63.525 176.880 63.560 ;
        RECT 175.950 62.990 176.280 63.390 ;
        RECT 176.705 63.160 177.235 63.525 ;
        RECT 177.425 63.160 177.700 64.010 ;
        RECT 177.870 63.160 178.060 64.520 ;
        RECT 178.230 64.535 178.400 65.200 ;
        RECT 178.570 64.780 178.740 65.540 ;
        RECT 178.975 64.780 179.490 65.190 ;
        RECT 178.230 64.345 178.980 64.535 ;
        RECT 179.150 63.970 179.490 64.780 ;
        RECT 179.660 64.450 180.870 65.540 ;
        RECT 178.260 63.800 179.490 63.970 ;
        RECT 178.240 62.990 178.750 63.525 ;
        RECT 178.970 63.195 179.215 63.800 ;
        RECT 179.660 63.740 180.180 64.280 ;
        RECT 180.350 63.910 180.870 64.450 ;
        RECT 181.045 64.400 181.380 65.370 ;
        RECT 181.550 64.400 181.720 65.540 ;
        RECT 181.890 65.200 183.920 65.370 ;
        RECT 179.660 62.990 180.870 63.740 ;
        RECT 181.045 63.730 181.215 64.400 ;
        RECT 181.890 64.230 182.060 65.200 ;
        RECT 181.385 63.900 181.640 64.230 ;
        RECT 181.865 63.900 182.060 64.230 ;
        RECT 182.230 64.860 183.355 65.030 ;
        RECT 181.470 63.730 181.640 63.900 ;
        RECT 182.230 63.730 182.400 64.860 ;
        RECT 181.045 63.160 181.300 63.730 ;
        RECT 181.470 63.560 182.400 63.730 ;
        RECT 182.570 64.520 183.580 64.690 ;
        RECT 182.570 63.720 182.740 64.520 ;
        RECT 182.225 63.525 182.400 63.560 ;
        RECT 181.470 62.990 181.800 63.390 ;
        RECT 182.225 63.160 182.755 63.525 ;
        RECT 182.945 63.500 183.220 64.320 ;
        RECT 182.940 63.330 183.220 63.500 ;
        RECT 182.945 63.160 183.220 63.330 ;
        RECT 183.390 63.160 183.580 64.520 ;
        RECT 183.750 64.535 183.920 65.200 ;
        RECT 184.090 64.780 184.260 65.540 ;
        RECT 184.495 64.780 185.010 65.190 ;
        RECT 185.180 65.105 190.525 65.540 ;
        RECT 183.750 64.345 184.500 64.535 ;
        RECT 184.670 63.970 185.010 64.780 ;
        RECT 183.780 63.800 185.010 63.970 ;
        RECT 183.760 62.990 184.270 63.525 ;
        RECT 184.490 63.195 184.735 63.800 ;
        RECT 186.765 63.535 187.105 64.365 ;
        RECT 188.585 63.855 188.935 65.105 ;
        RECT 190.700 64.450 193.290 65.540 ;
        RECT 190.700 63.760 191.910 64.280 ;
        RECT 192.080 63.930 193.290 64.450 ;
        RECT 193.995 64.570 194.270 65.370 ;
        RECT 194.440 64.740 194.770 65.540 ;
        RECT 194.940 65.200 196.020 65.370 ;
        RECT 194.940 64.570 195.110 65.200 ;
        RECT 193.995 64.360 195.110 64.570 ;
        RECT 195.325 64.520 195.570 65.030 ;
        RECT 195.740 64.700 196.020 65.200 ;
        RECT 196.255 64.700 196.505 65.540 ;
        RECT 196.720 64.520 196.890 65.370 ;
        RECT 197.060 64.780 197.390 65.540 ;
        RECT 198.060 65.030 199.250 65.320 ;
        RECT 197.625 64.570 197.795 64.820 ;
        RECT 195.325 64.350 196.890 64.520 ;
        RECT 197.110 64.400 197.795 64.570 ;
        RECT 198.080 64.690 199.250 64.860 ;
        RECT 199.420 64.740 199.700 65.540 ;
        RECT 198.080 64.400 198.405 64.690 ;
        RECT 199.080 64.570 199.250 64.690 ;
        RECT 193.920 63.980 194.715 64.180 ;
        RECT 194.885 63.980 196.025 64.180 ;
        RECT 196.195 63.810 196.450 64.350 ;
        RECT 197.110 64.150 197.280 64.400 ;
        RECT 198.575 64.230 198.770 64.520 ;
        RECT 199.080 64.400 199.740 64.570 ;
        RECT 199.910 64.400 200.185 65.370 ;
        RECT 199.570 64.230 199.740 64.400 ;
        RECT 196.640 63.980 197.280 64.150 ;
        RECT 185.180 62.990 190.525 63.535 ;
        RECT 190.700 62.990 193.290 63.760 ;
        RECT 193.995 63.630 195.950 63.810 ;
        RECT 193.995 63.170 194.350 63.630 ;
        RECT 194.520 62.990 194.690 63.460 ;
        RECT 194.860 63.160 195.190 63.630 ;
        RECT 195.360 62.990 195.530 63.460 ;
        RECT 195.700 63.380 195.950 63.630 ;
        RECT 196.120 63.550 196.450 63.810 ;
        RECT 196.620 63.380 196.900 63.810 ;
        RECT 195.700 63.160 196.900 63.380 ;
        RECT 197.110 63.730 197.280 63.980 ;
        RECT 197.450 63.900 197.890 64.230 ;
        RECT 198.060 63.900 198.405 64.230 ;
        RECT 198.575 63.900 199.400 64.230 ;
        RECT 199.570 63.900 199.845 64.230 ;
        RECT 199.570 63.730 199.740 63.900 ;
        RECT 197.110 63.350 197.375 63.730 ;
        RECT 197.625 62.990 197.795 63.730 ;
        RECT 198.075 63.560 199.740 63.730 ;
        RECT 200.015 63.665 200.185 64.400 ;
        RECT 200.820 64.375 201.110 65.540 ;
        RECT 201.280 64.400 201.620 65.370 ;
        RECT 201.790 64.400 201.960 65.540 ;
        RECT 202.230 64.740 202.480 65.540 ;
        RECT 203.125 64.570 203.455 65.370 ;
        RECT 203.755 64.740 204.085 65.540 ;
        RECT 204.255 64.570 204.585 65.370 ;
        RECT 202.150 64.400 204.585 64.570 ;
        RECT 204.960 64.450 206.630 65.540 ;
        RECT 201.280 63.790 201.455 64.400 ;
        RECT 202.150 64.150 202.320 64.400 ;
        RECT 201.625 63.980 202.320 64.150 ;
        RECT 202.495 63.980 202.915 64.180 ;
        RECT 203.085 63.980 203.415 64.180 ;
        RECT 203.585 63.980 203.915 64.180 ;
        RECT 198.075 63.210 198.330 63.560 ;
        RECT 198.500 62.990 198.830 63.390 ;
        RECT 199.000 63.210 199.170 63.560 ;
        RECT 199.340 62.990 199.720 63.390 ;
        RECT 199.910 63.320 200.185 63.665 ;
        RECT 200.820 62.990 201.110 63.715 ;
        RECT 201.280 63.160 201.620 63.790 ;
        RECT 201.790 62.990 202.040 63.790 ;
        RECT 202.230 63.640 203.455 63.810 ;
        RECT 202.230 63.160 202.560 63.640 ;
        RECT 202.730 62.990 202.955 63.450 ;
        RECT 203.125 63.160 203.455 63.640 ;
        RECT 204.085 63.770 204.255 64.400 ;
        RECT 204.440 63.980 204.790 64.230 ;
        RECT 204.085 63.160 204.585 63.770 ;
        RECT 204.960 63.760 205.710 64.280 ;
        RECT 205.880 63.930 206.630 64.450 ;
        RECT 207.465 64.570 207.795 65.370 ;
        RECT 207.965 64.740 208.295 65.540 ;
        RECT 208.595 64.570 208.925 65.370 ;
        RECT 209.570 64.740 209.820 65.540 ;
        RECT 207.465 64.400 209.900 64.570 ;
        RECT 210.090 64.400 210.260 65.540 ;
        RECT 210.430 64.400 210.770 65.370 ;
        RECT 211.145 64.570 211.475 65.370 ;
        RECT 211.645 64.740 211.975 65.540 ;
        RECT 212.275 64.570 212.605 65.370 ;
        RECT 213.250 64.740 213.500 65.540 ;
        RECT 211.145 64.400 213.580 64.570 ;
        RECT 213.770 64.400 213.940 65.540 ;
        RECT 214.110 64.400 214.450 65.370 ;
        RECT 214.825 64.570 215.155 65.370 ;
        RECT 215.325 64.740 215.655 65.540 ;
        RECT 215.955 64.570 216.285 65.370 ;
        RECT 216.930 64.740 217.180 65.540 ;
        RECT 214.825 64.400 217.260 64.570 ;
        RECT 217.450 64.400 217.620 65.540 ;
        RECT 217.790 64.400 218.130 65.370 ;
        RECT 207.260 63.980 207.610 64.230 ;
        RECT 207.795 63.770 207.965 64.400 ;
        RECT 208.135 63.980 208.465 64.180 ;
        RECT 208.635 63.980 208.965 64.180 ;
        RECT 209.135 63.980 209.555 64.180 ;
        RECT 209.730 64.150 209.900 64.400 ;
        RECT 210.540 64.350 210.770 64.400 ;
        RECT 209.730 63.980 210.425 64.150 ;
        RECT 204.960 62.990 206.630 63.760 ;
        RECT 207.465 63.160 207.965 63.770 ;
        RECT 208.595 63.640 209.820 63.810 ;
        RECT 210.595 63.790 210.770 64.350 ;
        RECT 210.940 63.980 211.290 64.230 ;
        RECT 208.595 63.160 208.925 63.640 ;
        RECT 209.095 62.990 209.320 63.450 ;
        RECT 209.490 63.160 209.820 63.640 ;
        RECT 210.010 62.990 210.260 63.790 ;
        RECT 210.430 63.160 210.770 63.790 ;
        RECT 211.475 63.770 211.645 64.400 ;
        RECT 211.815 63.980 212.145 64.180 ;
        RECT 212.315 63.980 212.645 64.180 ;
        RECT 212.815 63.980 213.235 64.180 ;
        RECT 213.410 64.150 213.580 64.400 ;
        RECT 213.410 63.980 214.105 64.150 ;
        RECT 214.275 63.840 214.450 64.400 ;
        RECT 214.620 63.980 214.970 64.230 ;
        RECT 211.145 63.160 211.645 63.770 ;
        RECT 212.275 63.640 213.500 63.810 ;
        RECT 214.220 63.790 214.450 63.840 ;
        RECT 212.275 63.160 212.605 63.640 ;
        RECT 212.775 62.990 213.000 63.450 ;
        RECT 213.170 63.160 213.500 63.640 ;
        RECT 213.690 62.990 213.940 63.790 ;
        RECT 214.110 63.160 214.450 63.790 ;
        RECT 215.155 63.770 215.325 64.400 ;
        RECT 215.495 63.980 215.825 64.180 ;
        RECT 215.995 63.980 216.325 64.180 ;
        RECT 216.495 63.980 216.915 64.180 ;
        RECT 217.090 64.150 217.260 64.400 ;
        RECT 217.090 63.980 217.785 64.150 ;
        RECT 217.955 63.840 218.130 64.400 ;
        RECT 214.825 63.160 215.325 63.770 ;
        RECT 215.955 63.640 217.180 63.810 ;
        RECT 217.900 63.790 218.130 63.840 ;
        RECT 215.955 63.160 216.285 63.640 ;
        RECT 216.455 62.990 216.680 63.450 ;
        RECT 216.850 63.160 217.180 63.640 ;
        RECT 217.370 62.990 217.620 63.790 ;
        RECT 217.790 63.160 218.130 63.790 ;
        RECT 218.300 64.400 218.685 65.360 ;
        RECT 218.900 64.740 219.190 65.540 ;
        RECT 219.360 65.200 220.725 65.370 ;
        RECT 219.360 64.570 219.530 65.200 ;
        RECT 218.855 64.400 219.530 64.570 ;
        RECT 218.300 63.730 218.475 64.400 ;
        RECT 218.855 64.230 219.025 64.400 ;
        RECT 219.700 64.230 220.025 65.030 ;
        RECT 220.395 64.990 220.725 65.200 ;
        RECT 220.395 64.740 221.350 64.990 ;
        RECT 218.660 63.980 219.025 64.230 ;
        RECT 219.220 63.980 219.470 64.230 ;
        RECT 218.660 63.900 218.850 63.980 ;
        RECT 219.220 63.900 219.390 63.980 ;
        RECT 219.680 63.900 220.025 64.230 ;
        RECT 220.195 63.900 220.470 64.565 ;
        RECT 220.655 63.900 221.010 64.565 ;
        RECT 221.180 63.730 221.350 64.740 ;
        RECT 221.520 64.400 221.810 65.540 ;
        RECT 221.980 64.450 225.490 65.540 ;
        RECT 221.535 63.900 221.810 64.230 ;
        RECT 218.300 63.160 218.810 63.730 ;
        RECT 219.355 63.560 220.755 63.730 ;
        RECT 218.980 62.990 219.150 63.550 ;
        RECT 219.355 63.160 219.685 63.560 ;
        RECT 219.860 62.990 220.190 63.390 ;
        RECT 220.425 63.370 220.755 63.560 ;
        RECT 220.925 63.540 221.350 63.730 ;
        RECT 221.980 63.760 223.630 64.280 ;
        RECT 223.800 63.930 225.490 64.450 ;
        RECT 226.580 64.375 226.870 65.540 ;
        RECT 227.040 65.105 232.385 65.540 ;
        RECT 232.560 65.105 237.905 65.540 ;
        RECT 221.520 63.370 221.810 63.640 ;
        RECT 220.425 63.160 221.810 63.370 ;
        RECT 221.980 62.990 225.490 63.760 ;
        RECT 226.580 62.990 226.870 63.715 ;
        RECT 228.625 63.535 228.965 64.365 ;
        RECT 230.445 63.855 230.795 65.105 ;
        RECT 234.145 63.535 234.485 64.365 ;
        RECT 235.965 63.855 236.315 65.105 ;
        RECT 238.080 64.450 240.670 65.540 ;
        RECT 238.080 63.760 239.290 64.280 ;
        RECT 239.460 63.930 240.670 64.450 ;
        RECT 241.350 64.525 241.605 65.365 ;
        RECT 241.780 64.720 242.110 65.540 ;
        RECT 242.350 64.550 242.560 65.365 ;
        RECT 227.040 62.990 232.385 63.535 ;
        RECT 232.560 62.990 237.905 63.535 ;
        RECT 238.080 62.990 240.670 63.760 ;
        RECT 241.350 63.160 241.680 64.525 ;
        RECT 241.910 64.370 242.560 64.550 ;
        RECT 241.910 63.730 242.130 64.370 ;
        RECT 242.730 64.195 242.935 65.370 ;
        RECT 242.505 63.955 242.935 64.195 ;
        RECT 243.105 63.955 243.435 65.370 ;
        RECT 243.615 63.900 243.895 65.370 ;
        RECT 244.075 64.570 244.360 65.365 ;
        RECT 244.540 64.740 244.755 65.540 ;
        RECT 244.935 64.570 245.205 65.365 ;
        RECT 245.440 65.105 250.785 65.540 ;
        RECT 244.075 64.400 245.205 64.570 ;
        RECT 244.120 63.900 244.505 64.230 ;
        RECT 244.725 63.930 245.225 64.195 ;
        RECT 244.200 63.750 244.505 63.900 ;
        RECT 241.910 63.560 244.020 63.730 ;
        RECT 241.910 63.555 243.130 63.560 ;
        RECT 241.850 62.990 242.525 63.375 ;
        RECT 242.800 63.165 243.130 63.555 ;
        RECT 243.300 62.990 243.645 63.390 ;
        RECT 243.815 63.165 244.020 63.560 ;
        RECT 244.200 63.190 244.755 63.750 ;
        RECT 244.930 62.990 245.170 63.665 ;
        RECT 247.025 63.535 247.365 64.365 ;
        RECT 248.845 63.855 249.195 65.105 ;
        RECT 250.960 64.450 252.170 65.540 ;
        RECT 250.960 63.740 251.480 64.280 ;
        RECT 251.650 63.910 252.170 64.450 ;
        RECT 252.340 64.375 252.630 65.540 ;
        RECT 252.800 64.450 256.310 65.540 ;
        RECT 252.800 63.760 254.450 64.280 ;
        RECT 254.620 63.930 256.310 64.450 ;
        RECT 256.940 63.935 257.220 65.370 ;
        RECT 257.390 64.765 258.100 65.540 ;
        RECT 258.270 64.595 258.600 65.370 ;
        RECT 257.450 64.380 258.600 64.595 ;
        RECT 245.440 62.990 250.785 63.535 ;
        RECT 250.960 62.990 252.170 63.740 ;
        RECT 252.340 62.990 252.630 63.715 ;
        RECT 252.800 62.990 256.310 63.760 ;
        RECT 256.940 63.160 257.280 63.935 ;
        RECT 257.450 63.810 257.735 64.380 ;
        RECT 257.920 63.980 258.390 64.210 ;
        RECT 258.795 64.180 259.010 65.295 ;
        RECT 259.190 64.820 259.520 65.540 ;
        RECT 259.700 65.105 265.045 65.540 ;
        RECT 265.220 65.105 270.565 65.540 ;
        RECT 259.300 64.180 259.530 64.520 ;
        RECT 258.560 64.000 259.010 64.180 ;
        RECT 258.560 63.980 258.890 64.000 ;
        RECT 259.200 63.980 259.530 64.180 ;
        RECT 257.450 63.620 258.160 63.810 ;
        RECT 257.860 63.480 258.160 63.620 ;
        RECT 258.350 63.620 259.530 63.810 ;
        RECT 258.350 63.540 258.680 63.620 ;
        RECT 257.860 63.470 258.175 63.480 ;
        RECT 257.860 63.460 258.185 63.470 ;
        RECT 257.860 63.455 258.195 63.460 ;
        RECT 257.450 62.990 257.620 63.450 ;
        RECT 257.860 63.445 258.200 63.455 ;
        RECT 257.860 63.440 258.205 63.445 ;
        RECT 257.860 63.430 258.210 63.440 ;
        RECT 257.860 63.425 258.215 63.430 ;
        RECT 257.860 63.160 258.220 63.425 ;
        RECT 258.850 62.990 259.020 63.450 ;
        RECT 259.190 63.160 259.530 63.620 ;
        RECT 261.285 63.535 261.625 64.365 ;
        RECT 263.105 63.855 263.455 65.105 ;
        RECT 266.805 63.535 267.145 64.365 ;
        RECT 268.625 63.855 268.975 65.105 ;
        RECT 270.740 64.450 271.950 65.540 ;
        RECT 272.120 65.035 272.750 65.540 ;
        RECT 270.740 63.740 271.260 64.280 ;
        RECT 271.430 63.910 271.950 64.450 ;
        RECT 272.135 64.500 272.390 64.865 ;
        RECT 272.560 64.860 272.750 65.035 ;
        RECT 272.930 65.030 273.405 65.370 ;
        RECT 272.560 64.670 272.890 64.860 ;
        RECT 273.115 64.500 273.365 64.795 ;
        RECT 273.590 64.695 273.805 65.540 ;
        RECT 274.005 64.700 274.280 65.370 ;
        RECT 272.135 64.330 273.925 64.500 ;
        RECT 274.110 64.350 274.280 64.700 ;
        RECT 274.450 64.530 274.710 65.540 ;
        RECT 274.880 64.450 277.470 65.540 ;
        RECT 259.700 62.990 265.045 63.535 ;
        RECT 265.220 62.990 270.565 63.535 ;
        RECT 270.740 62.990 271.950 63.740 ;
        RECT 272.120 63.670 272.505 64.150 ;
        RECT 272.675 63.475 272.930 64.330 ;
        RECT 272.140 63.210 272.930 63.475 ;
        RECT 273.100 63.655 273.510 64.150 ;
        RECT 273.695 63.900 273.925 64.330 ;
        RECT 274.095 63.830 274.710 64.350 ;
        RECT 273.100 63.210 273.330 63.655 ;
        RECT 274.095 63.620 274.265 63.830 ;
        RECT 274.880 63.760 276.090 64.280 ;
        RECT 276.260 63.930 277.470 64.450 ;
        RECT 278.100 64.375 278.390 65.540 ;
        RECT 278.560 64.450 280.230 65.540 ;
        RECT 280.405 64.870 280.660 65.370 ;
        RECT 280.830 65.040 281.160 65.540 ;
        RECT 280.405 64.700 281.155 64.870 ;
        RECT 278.560 63.760 279.310 64.280 ;
        RECT 279.480 63.930 280.230 64.450 ;
        RECT 280.405 63.880 280.755 64.530 ;
        RECT 273.510 62.990 273.840 63.485 ;
        RECT 274.015 63.160 274.265 63.620 ;
        RECT 274.435 62.990 274.710 63.650 ;
        RECT 274.880 62.990 277.470 63.760 ;
        RECT 278.100 62.990 278.390 63.715 ;
        RECT 278.560 62.990 280.230 63.760 ;
        RECT 280.925 63.710 281.155 64.700 ;
        RECT 280.405 63.540 281.155 63.710 ;
        RECT 280.405 63.250 280.660 63.540 ;
        RECT 280.830 62.990 281.160 63.370 ;
        RECT 281.330 63.250 281.500 65.370 ;
        RECT 281.670 64.570 281.995 65.355 ;
        RECT 282.165 65.080 282.415 65.540 ;
        RECT 282.585 65.040 282.835 65.370 ;
        RECT 283.050 65.040 283.730 65.370 ;
        RECT 282.585 64.910 282.755 65.040 ;
        RECT 282.360 64.740 282.755 64.910 ;
        RECT 281.730 63.520 282.190 64.570 ;
        RECT 282.360 63.380 282.530 64.740 ;
        RECT 282.925 64.480 283.390 64.870 ;
        RECT 282.700 63.670 283.050 64.290 ;
        RECT 283.220 63.890 283.390 64.480 ;
        RECT 283.560 64.260 283.730 65.040 ;
        RECT 283.900 64.940 284.070 65.280 ;
        RECT 284.305 65.110 284.635 65.540 ;
        RECT 284.805 64.940 284.975 65.280 ;
        RECT 285.270 65.080 285.640 65.540 ;
        RECT 283.900 64.770 284.975 64.940 ;
        RECT 285.810 64.910 285.980 65.370 ;
        RECT 286.215 65.030 287.085 65.370 ;
        RECT 287.255 65.080 287.505 65.540 ;
        RECT 285.420 64.740 285.980 64.910 ;
        RECT 285.420 64.600 285.590 64.740 ;
        RECT 284.090 64.430 285.590 64.600 ;
        RECT 286.285 64.570 286.745 64.860 ;
        RECT 283.560 64.090 285.250 64.260 ;
        RECT 283.220 63.670 283.575 63.890 ;
        RECT 283.745 63.380 283.915 64.090 ;
        RECT 284.120 63.670 284.910 63.920 ;
        RECT 285.080 63.910 285.250 64.090 ;
        RECT 285.420 63.740 285.590 64.430 ;
        RECT 281.860 62.990 282.190 63.350 ;
        RECT 282.360 63.210 282.855 63.380 ;
        RECT 283.060 63.210 283.915 63.380 ;
        RECT 284.790 62.990 285.120 63.450 ;
        RECT 285.330 63.350 285.590 63.740 ;
        RECT 285.780 64.560 286.745 64.570 ;
        RECT 286.915 64.650 287.085 65.030 ;
        RECT 287.675 64.990 287.845 65.280 ;
        RECT 288.025 65.160 288.355 65.540 ;
        RECT 287.675 64.820 288.475 64.990 ;
        RECT 285.780 64.400 286.455 64.560 ;
        RECT 286.915 64.480 288.135 64.650 ;
        RECT 285.780 63.610 285.990 64.400 ;
        RECT 286.915 64.390 287.085 64.480 ;
        RECT 286.160 63.610 286.510 64.230 ;
        RECT 286.680 64.220 287.085 64.390 ;
        RECT 286.680 63.440 286.850 64.220 ;
        RECT 287.020 63.770 287.240 64.050 ;
        RECT 287.420 63.940 287.960 64.310 ;
        RECT 288.305 64.230 288.475 64.820 ;
        RECT 288.695 64.400 289.000 65.540 ;
        RECT 289.170 64.350 289.425 65.230 ;
        RECT 289.600 64.450 293.110 65.540 ;
        RECT 294.205 64.870 294.460 65.370 ;
        RECT 294.630 65.040 294.960 65.540 ;
        RECT 294.205 64.700 294.955 64.870 ;
        RECT 288.305 64.200 289.045 64.230 ;
        RECT 287.020 63.600 287.550 63.770 ;
        RECT 285.330 63.180 285.680 63.350 ;
        RECT 285.900 63.160 286.850 63.440 ;
        RECT 287.020 62.990 287.210 63.430 ;
        RECT 287.380 63.370 287.550 63.600 ;
        RECT 287.720 63.540 287.960 63.940 ;
        RECT 288.130 63.900 289.045 64.200 ;
        RECT 288.130 63.725 288.455 63.900 ;
        RECT 288.130 63.370 288.450 63.725 ;
        RECT 289.215 63.700 289.425 64.350 ;
        RECT 287.380 63.200 288.450 63.370 ;
        RECT 288.695 62.990 289.000 63.450 ;
        RECT 289.170 63.170 289.425 63.700 ;
        RECT 289.600 63.760 291.250 64.280 ;
        RECT 291.420 63.930 293.110 64.450 ;
        RECT 294.205 63.880 294.555 64.530 ;
        RECT 289.600 62.990 293.110 63.760 ;
        RECT 294.725 63.710 294.955 64.700 ;
        RECT 294.205 63.540 294.955 63.710 ;
        RECT 294.205 63.250 294.460 63.540 ;
        RECT 294.630 62.990 294.960 63.370 ;
        RECT 295.130 63.250 295.300 65.370 ;
        RECT 295.470 64.570 295.795 65.355 ;
        RECT 295.965 65.080 296.215 65.540 ;
        RECT 296.385 65.040 296.635 65.370 ;
        RECT 296.850 65.040 297.530 65.370 ;
        RECT 296.385 64.910 296.555 65.040 ;
        RECT 296.160 64.740 296.555 64.910 ;
        RECT 295.530 63.520 295.990 64.570 ;
        RECT 296.160 63.380 296.330 64.740 ;
        RECT 296.725 64.480 297.190 64.870 ;
        RECT 296.500 63.670 296.850 64.290 ;
        RECT 297.020 63.890 297.190 64.480 ;
        RECT 297.360 64.260 297.530 65.040 ;
        RECT 297.700 64.940 297.870 65.280 ;
        RECT 298.105 65.110 298.435 65.540 ;
        RECT 298.605 64.940 298.775 65.280 ;
        RECT 299.070 65.080 299.440 65.540 ;
        RECT 297.700 64.770 298.775 64.940 ;
        RECT 299.610 64.910 299.780 65.370 ;
        RECT 300.015 65.030 300.885 65.370 ;
        RECT 301.055 65.080 301.305 65.540 ;
        RECT 299.220 64.740 299.780 64.910 ;
        RECT 299.220 64.600 299.390 64.740 ;
        RECT 297.890 64.430 299.390 64.600 ;
        RECT 300.085 64.570 300.545 64.860 ;
        RECT 297.360 64.090 299.050 64.260 ;
        RECT 297.020 63.670 297.375 63.890 ;
        RECT 297.545 63.380 297.715 64.090 ;
        RECT 297.920 63.670 298.710 63.920 ;
        RECT 298.880 63.910 299.050 64.090 ;
        RECT 299.220 63.740 299.390 64.430 ;
        RECT 295.660 62.990 295.990 63.350 ;
        RECT 296.160 63.210 296.655 63.380 ;
        RECT 296.860 63.210 297.715 63.380 ;
        RECT 298.590 62.990 298.920 63.450 ;
        RECT 299.130 63.350 299.390 63.740 ;
        RECT 299.580 64.560 300.545 64.570 ;
        RECT 300.715 64.650 300.885 65.030 ;
        RECT 301.475 64.990 301.645 65.280 ;
        RECT 301.825 65.160 302.155 65.540 ;
        RECT 301.475 64.820 302.275 64.990 ;
        RECT 299.580 64.400 300.255 64.560 ;
        RECT 300.715 64.480 301.935 64.650 ;
        RECT 299.580 63.610 299.790 64.400 ;
        RECT 300.715 64.390 300.885 64.480 ;
        RECT 299.960 63.610 300.310 64.230 ;
        RECT 300.480 64.220 300.885 64.390 ;
        RECT 300.480 63.440 300.650 64.220 ;
        RECT 300.820 63.770 301.040 64.050 ;
        RECT 301.220 63.940 301.760 64.310 ;
        RECT 302.105 64.230 302.275 64.820 ;
        RECT 302.495 64.400 302.800 65.540 ;
        RECT 302.970 64.350 303.220 65.230 ;
        RECT 303.390 64.400 303.640 65.540 ;
        RECT 303.860 64.375 304.150 65.540 ;
        RECT 304.325 64.400 304.660 65.370 ;
        RECT 304.830 64.400 305.000 65.540 ;
        RECT 305.170 65.200 307.200 65.370 ;
        RECT 302.105 64.200 302.845 64.230 ;
        RECT 300.820 63.600 301.350 63.770 ;
        RECT 299.130 63.180 299.480 63.350 ;
        RECT 299.700 63.160 300.650 63.440 ;
        RECT 300.820 62.990 301.010 63.430 ;
        RECT 301.180 63.370 301.350 63.600 ;
        RECT 301.520 63.540 301.760 63.940 ;
        RECT 301.930 63.900 302.845 64.200 ;
        RECT 301.930 63.725 302.255 63.900 ;
        RECT 301.930 63.370 302.250 63.725 ;
        RECT 303.015 63.700 303.220 64.350 ;
        RECT 301.180 63.200 302.250 63.370 ;
        RECT 302.495 62.990 302.800 63.450 ;
        RECT 302.970 63.170 303.220 63.700 ;
        RECT 303.390 62.990 303.640 63.745 ;
        RECT 304.325 63.730 304.495 64.400 ;
        RECT 305.170 64.230 305.340 65.200 ;
        RECT 304.665 63.900 304.920 64.230 ;
        RECT 305.145 63.900 305.340 64.230 ;
        RECT 305.510 64.860 306.635 65.030 ;
        RECT 304.750 63.730 304.920 63.900 ;
        RECT 305.510 63.730 305.680 64.860 ;
        RECT 303.860 62.990 304.150 63.715 ;
        RECT 304.325 63.160 304.580 63.730 ;
        RECT 304.750 63.560 305.680 63.730 ;
        RECT 305.850 64.520 306.860 64.690 ;
        RECT 305.850 63.720 306.020 64.520 ;
        RECT 306.225 64.180 306.500 64.320 ;
        RECT 306.220 64.010 306.500 64.180 ;
        RECT 305.505 63.525 305.680 63.560 ;
        RECT 304.750 62.990 305.080 63.390 ;
        RECT 305.505 63.160 306.035 63.525 ;
        RECT 306.225 63.160 306.500 64.010 ;
        RECT 306.670 63.160 306.860 64.520 ;
        RECT 307.030 64.535 307.200 65.200 ;
        RECT 307.370 64.780 307.540 65.540 ;
        RECT 307.775 64.780 308.290 65.190 ;
        RECT 307.030 64.345 307.780 64.535 ;
        RECT 307.950 63.970 308.290 64.780 ;
        RECT 308.460 64.450 309.670 65.540 ;
        RECT 307.060 63.800 308.290 63.970 ;
        RECT 307.040 62.990 307.550 63.525 ;
        RECT 307.770 63.195 308.015 63.800 ;
        RECT 308.460 63.740 308.980 64.280 ;
        RECT 309.150 63.910 309.670 64.450 ;
        RECT 309.840 64.450 311.050 65.540 ;
        RECT 309.840 63.910 310.360 64.450 ;
        RECT 310.530 63.740 311.050 64.280 ;
        RECT 308.460 62.990 309.670 63.740 ;
        RECT 309.840 62.990 311.050 63.740 ;
        RECT 162.095 62.820 311.135 62.990 ;
        RECT 162.180 62.070 163.390 62.820 ;
        RECT 162.180 61.530 162.700 62.070 ;
        RECT 163.565 61.980 163.825 62.820 ;
        RECT 164.000 62.075 164.255 62.650 ;
        RECT 164.425 62.440 164.755 62.820 ;
        RECT 164.970 62.270 165.140 62.650 ;
        RECT 164.425 62.100 165.140 62.270 ;
        RECT 162.870 61.360 163.390 61.900 ;
        RECT 162.180 60.270 163.390 61.360 ;
        RECT 163.565 60.270 163.825 61.420 ;
        RECT 164.000 61.345 164.170 62.075 ;
        RECT 164.425 61.910 164.595 62.100 ;
        RECT 165.400 62.050 167.990 62.820 ;
        RECT 168.210 62.065 168.460 62.820 ;
        RECT 168.630 62.110 168.880 62.640 ;
        RECT 169.050 62.360 169.355 62.820 ;
        RECT 169.600 62.440 170.670 62.610 ;
        RECT 164.340 61.580 164.595 61.910 ;
        RECT 164.425 61.370 164.595 61.580 ;
        RECT 164.875 61.550 165.230 61.920 ;
        RECT 165.400 61.530 166.610 62.050 ;
        RECT 164.000 60.440 164.255 61.345 ;
        RECT 164.425 61.200 165.140 61.370 ;
        RECT 166.780 61.360 167.990 61.880 ;
        RECT 168.630 61.460 168.835 62.110 ;
        RECT 169.600 62.085 169.920 62.440 ;
        RECT 169.595 61.910 169.920 62.085 ;
        RECT 169.005 61.610 169.920 61.910 ;
        RECT 170.090 61.870 170.330 62.270 ;
        RECT 170.500 62.210 170.670 62.440 ;
        RECT 170.840 62.380 171.030 62.820 ;
        RECT 171.200 62.370 172.150 62.650 ;
        RECT 172.370 62.460 172.720 62.630 ;
        RECT 170.500 62.040 171.030 62.210 ;
        RECT 169.005 61.580 169.745 61.610 ;
        RECT 164.425 60.270 164.755 61.030 ;
        RECT 164.970 60.440 165.140 61.200 ;
        RECT 165.400 60.270 167.990 61.360 ;
        RECT 168.210 60.270 168.460 61.410 ;
        RECT 168.630 60.580 168.880 61.460 ;
        RECT 169.050 60.270 169.355 61.410 ;
        RECT 169.575 60.990 169.745 61.580 ;
        RECT 170.090 61.500 170.630 61.870 ;
        RECT 170.810 61.760 171.030 62.040 ;
        RECT 171.200 61.590 171.370 62.370 ;
        RECT 170.965 61.420 171.370 61.590 ;
        RECT 171.540 61.580 171.890 62.200 ;
        RECT 170.965 61.330 171.135 61.420 ;
        RECT 172.060 61.410 172.270 62.200 ;
        RECT 169.915 61.160 171.135 61.330 ;
        RECT 171.595 61.250 172.270 61.410 ;
        RECT 169.575 60.820 170.375 60.990 ;
        RECT 169.695 60.270 170.025 60.650 ;
        RECT 170.205 60.530 170.375 60.820 ;
        RECT 170.965 60.780 171.135 61.160 ;
        RECT 171.305 61.240 172.270 61.250 ;
        RECT 172.460 62.070 172.720 62.460 ;
        RECT 172.930 62.360 173.260 62.820 ;
        RECT 174.135 62.430 174.990 62.600 ;
        RECT 175.195 62.430 175.690 62.600 ;
        RECT 175.860 62.460 176.190 62.820 ;
        RECT 172.460 61.380 172.630 62.070 ;
        RECT 172.800 61.720 172.970 61.900 ;
        RECT 173.140 61.890 173.930 62.140 ;
        RECT 174.135 61.720 174.305 62.430 ;
        RECT 174.475 61.920 174.830 62.140 ;
        RECT 172.800 61.550 174.490 61.720 ;
        RECT 171.305 60.950 171.765 61.240 ;
        RECT 172.460 61.210 173.960 61.380 ;
        RECT 172.460 61.070 172.630 61.210 ;
        RECT 172.070 60.900 172.630 61.070 ;
        RECT 170.545 60.270 170.795 60.730 ;
        RECT 170.965 60.440 171.835 60.780 ;
        RECT 172.070 60.440 172.240 60.900 ;
        RECT 173.075 60.870 174.150 61.040 ;
        RECT 172.410 60.270 172.780 60.730 ;
        RECT 173.075 60.530 173.245 60.870 ;
        RECT 173.415 60.270 173.745 60.700 ;
        RECT 173.980 60.530 174.150 60.870 ;
        RECT 174.320 60.770 174.490 61.550 ;
        RECT 174.660 61.330 174.830 61.920 ;
        RECT 175.000 61.520 175.350 62.140 ;
        RECT 174.660 60.940 175.125 61.330 ;
        RECT 175.520 61.070 175.690 62.430 ;
        RECT 175.860 61.240 176.320 62.290 ;
        RECT 175.295 60.900 175.690 61.070 ;
        RECT 175.295 60.770 175.465 60.900 ;
        RECT 174.320 60.440 175.000 60.770 ;
        RECT 175.215 60.440 175.465 60.770 ;
        RECT 175.635 60.270 175.885 60.730 ;
        RECT 176.055 60.455 176.380 61.240 ;
        RECT 176.550 60.440 176.720 62.560 ;
        RECT 176.890 62.440 177.220 62.820 ;
        RECT 177.390 62.270 177.645 62.560 ;
        RECT 176.895 62.100 177.645 62.270 ;
        RECT 176.895 61.110 177.125 62.100 ;
        RECT 177.820 62.020 178.110 62.820 ;
        RECT 178.280 62.360 178.830 62.650 ;
        RECT 179.000 62.360 179.250 62.820 ;
        RECT 177.295 61.280 177.645 61.930 ;
        RECT 176.895 60.940 177.645 61.110 ;
        RECT 176.890 60.270 177.220 60.770 ;
        RECT 177.390 60.440 177.645 60.940 ;
        RECT 177.820 60.270 178.110 61.410 ;
        RECT 178.280 60.990 178.530 62.360 ;
        RECT 179.880 62.190 180.210 62.550 ;
        RECT 178.820 62.000 180.210 62.190 ;
        RECT 180.580 62.050 184.090 62.820 ;
        RECT 184.790 62.420 185.120 62.820 ;
        RECT 185.290 62.250 185.460 62.520 ;
        RECT 185.630 62.420 185.960 62.820 ;
        RECT 186.130 62.250 186.385 62.520 ;
        RECT 178.820 61.910 178.990 62.000 ;
        RECT 178.700 61.580 178.990 61.910 ;
        RECT 179.160 61.580 179.490 61.830 ;
        RECT 179.720 61.580 180.410 61.830 ;
        RECT 178.820 61.330 178.990 61.580 ;
        RECT 178.820 61.160 179.760 61.330 ;
        RECT 178.280 60.440 178.730 60.990 ;
        RECT 178.920 60.270 179.250 60.990 ;
        RECT 179.460 60.610 179.760 61.160 ;
        RECT 180.095 61.140 180.410 61.580 ;
        RECT 180.580 61.530 182.230 62.050 ;
        RECT 182.400 61.360 184.090 61.880 ;
        RECT 179.930 60.270 180.210 60.940 ;
        RECT 180.580 60.270 184.090 61.360 ;
        RECT 184.720 61.240 184.990 62.250 ;
        RECT 185.160 62.080 186.385 62.250 ;
        RECT 185.160 61.410 185.330 62.080 ;
        RECT 186.560 62.070 187.770 62.820 ;
        RECT 187.940 62.095 188.230 62.820 ;
        RECT 188.860 62.440 189.190 62.820 ;
        RECT 188.415 62.270 188.690 62.410 ;
        RECT 189.360 62.270 189.570 62.440 ;
        RECT 188.415 62.080 189.570 62.270 ;
        RECT 189.740 62.270 190.070 62.650 ;
        RECT 190.260 62.440 190.590 62.820 ;
        RECT 185.500 61.580 185.880 61.910 ;
        RECT 186.050 61.580 186.385 61.910 ;
        RECT 185.160 61.240 185.475 61.410 ;
        RECT 184.725 60.270 185.040 61.070 ;
        RECT 185.305 60.625 185.475 61.240 ;
        RECT 185.645 60.900 185.880 61.580 ;
        RECT 186.560 61.530 187.080 62.070 ;
        RECT 189.740 62.065 190.590 62.270 ;
        RECT 186.050 60.625 186.385 61.410 ;
        RECT 187.250 61.360 187.770 61.900 ;
        RECT 188.410 61.455 188.670 61.910 ;
        RECT 188.925 61.505 189.510 61.880 ;
        RECT 185.305 60.455 186.385 60.625 ;
        RECT 186.560 60.270 187.770 61.360 ;
        RECT 187.940 60.270 188.230 61.435 ;
        RECT 188.415 60.270 188.740 61.255 ;
        RECT 188.925 61.120 189.130 61.505 ;
        RECT 189.680 61.290 190.090 61.895 ;
        RECT 190.260 61.575 190.590 62.065 ;
        RECT 190.260 61.120 190.430 61.575 ;
        RECT 188.920 60.950 189.130 61.120 ;
        RECT 188.925 60.920 189.130 60.950 ;
        RECT 189.310 60.900 190.430 61.120 ;
        RECT 189.310 60.440 189.570 60.900 ;
        RECT 189.740 60.270 190.590 60.720 ;
        RECT 190.760 60.440 191.005 62.650 ;
        RECT 191.190 62.020 191.430 62.820 ;
        RECT 192.550 62.315 192.880 62.820 ;
        RECT 193.050 62.250 193.290 62.625 ;
        RECT 193.570 62.490 193.740 62.635 ;
        RECT 193.570 62.295 193.970 62.490 ;
        RECT 194.330 62.325 194.730 62.820 ;
        RECT 192.605 61.800 192.905 62.140 ;
        RECT 192.600 61.630 192.905 61.800 ;
        RECT 192.605 61.290 192.905 61.630 ;
        RECT 193.075 62.100 193.290 62.250 ;
        RECT 193.075 61.770 193.630 62.100 ;
        RECT 193.800 61.960 193.970 62.295 ;
        RECT 194.900 62.130 195.135 62.650 ;
        RECT 195.320 62.185 195.590 62.820 ;
        RECT 191.190 60.270 191.445 61.270 ;
        RECT 193.075 61.120 193.310 61.770 ;
        RECT 193.800 61.600 194.790 61.960 ;
        RECT 192.630 60.890 193.310 61.120 ;
        RECT 193.500 61.580 194.790 61.600 ;
        RECT 193.500 61.430 194.360 61.580 ;
        RECT 192.630 60.460 192.800 60.890 ;
        RECT 192.970 60.270 193.300 60.720 ;
        RECT 193.500 60.485 193.785 61.430 ;
        RECT 194.960 61.325 195.135 62.130 ;
        RECT 193.960 60.950 194.655 61.260 ;
        RECT 193.965 60.270 194.650 60.740 ;
        RECT 194.830 60.540 195.135 61.325 ;
        RECT 196.220 62.020 196.560 62.650 ;
        RECT 196.850 62.360 197.020 62.820 ;
        RECT 197.290 62.190 197.620 62.635 ;
        RECT 196.220 61.450 196.490 62.020 ;
        RECT 196.870 62.000 197.620 62.190 ;
        RECT 197.790 62.170 197.960 62.490 ;
        RECT 198.185 62.360 198.515 62.820 ;
        RECT 198.715 62.170 199.045 62.650 ;
        RECT 199.260 62.360 199.590 62.820 ;
        RECT 199.760 62.170 200.090 62.650 ;
        RECT 197.790 62.000 200.090 62.170 ;
        RECT 200.560 62.190 200.890 62.550 ;
        RECT 201.510 62.360 201.760 62.820 ;
        RECT 201.930 62.360 202.490 62.650 ;
        RECT 200.560 62.000 201.950 62.190 ;
        RECT 196.870 61.830 197.240 62.000 ;
        RECT 201.780 61.910 201.950 62.000 ;
        RECT 196.660 61.620 197.240 61.830 ;
        RECT 197.410 61.620 197.830 61.830 ;
        RECT 196.980 61.450 197.240 61.620 ;
        RECT 195.320 60.270 195.590 61.225 ;
        RECT 196.220 60.440 196.745 61.450 ;
        RECT 196.980 61.160 197.730 61.450 ;
        RECT 196.980 60.270 197.310 60.990 ;
        RECT 197.480 60.440 197.730 61.160 ;
        RECT 198.000 60.515 198.330 61.830 ;
        RECT 198.540 60.515 198.870 61.830 ;
        RECT 199.040 60.515 199.410 61.830 ;
        RECT 199.620 61.580 200.130 61.830 ;
        RECT 200.375 61.580 201.050 61.830 ;
        RECT 201.270 61.580 201.610 61.830 ;
        RECT 201.780 61.580 202.070 61.910 ;
        RECT 199.740 60.270 200.070 61.390 ;
        RECT 200.375 61.220 200.640 61.580 ;
        RECT 201.780 61.330 201.950 61.580 ;
        RECT 201.010 61.160 201.950 61.330 ;
        RECT 200.560 60.270 200.840 60.940 ;
        RECT 201.010 60.610 201.310 61.160 ;
        RECT 202.240 60.990 202.490 62.360 ;
        RECT 202.660 62.050 206.170 62.820 ;
        RECT 202.660 61.530 204.310 62.050 ;
        RECT 207.260 62.020 207.600 62.650 ;
        RECT 207.890 62.360 208.060 62.820 ;
        RECT 208.330 62.190 208.660 62.635 ;
        RECT 204.480 61.360 206.170 61.880 ;
        RECT 201.510 60.270 201.840 60.990 ;
        RECT 202.030 60.440 202.490 60.990 ;
        RECT 202.660 60.270 206.170 61.360 ;
        RECT 207.260 61.450 207.530 62.020 ;
        RECT 207.910 62.000 208.660 62.190 ;
        RECT 208.830 62.170 209.000 62.490 ;
        RECT 209.225 62.360 209.555 62.820 ;
        RECT 209.755 62.170 210.085 62.650 ;
        RECT 210.300 62.360 210.630 62.820 ;
        RECT 210.800 62.170 211.130 62.650 ;
        RECT 208.830 62.000 211.130 62.170 ;
        RECT 211.400 62.360 211.960 62.650 ;
        RECT 212.130 62.360 212.380 62.820 ;
        RECT 207.910 61.830 208.280 62.000 ;
        RECT 207.700 61.620 208.280 61.830 ;
        RECT 208.450 61.620 208.870 61.830 ;
        RECT 208.020 61.450 208.280 61.620 ;
        RECT 207.260 60.440 207.785 61.450 ;
        RECT 208.020 61.160 208.770 61.450 ;
        RECT 208.020 60.270 208.350 60.990 ;
        RECT 208.520 60.440 208.770 61.160 ;
        RECT 209.040 60.515 209.370 61.830 ;
        RECT 209.580 60.515 209.910 61.830 ;
        RECT 210.080 60.515 210.450 61.830 ;
        RECT 210.660 61.580 211.170 61.830 ;
        RECT 210.780 60.270 211.110 61.390 ;
        RECT 211.400 60.990 211.650 62.360 ;
        RECT 213.000 62.190 213.330 62.550 ;
        RECT 211.940 62.000 213.330 62.190 ;
        RECT 213.700 62.095 213.990 62.820 ;
        RECT 214.160 62.020 214.500 62.650 ;
        RECT 214.790 62.360 214.960 62.820 ;
        RECT 215.230 62.190 215.560 62.635 ;
        RECT 211.940 61.910 212.110 62.000 ;
        RECT 211.820 61.580 212.110 61.910 ;
        RECT 212.280 61.580 212.620 61.830 ;
        RECT 212.840 61.580 213.515 61.830 ;
        RECT 211.940 61.330 212.110 61.580 ;
        RECT 211.940 61.160 212.880 61.330 ;
        RECT 213.250 61.220 213.515 61.580 ;
        RECT 214.160 61.450 214.430 62.020 ;
        RECT 214.810 62.000 215.560 62.190 ;
        RECT 215.730 62.170 215.900 62.490 ;
        RECT 216.125 62.360 216.455 62.820 ;
        RECT 216.655 62.170 216.985 62.650 ;
        RECT 217.200 62.360 217.530 62.820 ;
        RECT 217.700 62.170 218.030 62.650 ;
        RECT 215.730 62.000 218.030 62.170 ;
        RECT 218.300 62.050 220.890 62.820 ;
        RECT 221.635 62.190 221.920 62.650 ;
        RECT 222.090 62.360 222.360 62.820 ;
        RECT 214.810 61.830 215.180 62.000 ;
        RECT 214.600 61.620 215.180 61.830 ;
        RECT 215.350 61.620 215.770 61.830 ;
        RECT 214.920 61.450 215.180 61.620 ;
        RECT 211.400 60.440 211.860 60.990 ;
        RECT 212.050 60.270 212.380 60.990 ;
        RECT 212.580 60.610 212.880 61.160 ;
        RECT 213.050 60.270 213.330 60.940 ;
        RECT 213.700 60.270 213.990 61.435 ;
        RECT 214.160 60.440 214.685 61.450 ;
        RECT 214.920 61.160 215.670 61.450 ;
        RECT 214.920 60.270 215.250 60.990 ;
        RECT 215.420 60.440 215.670 61.160 ;
        RECT 215.940 60.515 216.270 61.830 ;
        RECT 216.480 60.515 216.810 61.830 ;
        RECT 216.980 60.515 217.350 61.830 ;
        RECT 217.560 61.580 218.070 61.830 ;
        RECT 218.300 61.530 219.510 62.050 ;
        RECT 221.635 62.020 222.590 62.190 ;
        RECT 217.680 60.270 218.010 61.390 ;
        RECT 219.680 61.360 220.890 61.880 ;
        RECT 218.300 60.270 220.890 61.360 ;
        RECT 221.520 61.290 222.210 61.850 ;
        RECT 222.380 61.120 222.590 62.020 ;
        RECT 221.635 60.900 222.590 61.120 ;
        RECT 222.760 61.850 223.160 62.650 ;
        RECT 223.350 62.190 223.630 62.650 ;
        RECT 224.150 62.360 224.475 62.820 ;
        RECT 223.350 62.020 224.475 62.190 ;
        RECT 224.645 62.080 225.030 62.650 ;
        RECT 224.025 61.910 224.475 62.020 ;
        RECT 222.760 61.290 223.855 61.850 ;
        RECT 224.025 61.580 224.580 61.910 ;
        RECT 221.635 60.440 221.920 60.900 ;
        RECT 222.090 60.270 222.360 60.730 ;
        RECT 222.760 60.440 223.160 61.290 ;
        RECT 224.025 61.120 224.475 61.580 ;
        RECT 224.750 61.410 225.030 62.080 ;
        RECT 223.350 60.900 224.475 61.120 ;
        RECT 223.350 60.440 223.630 60.900 ;
        RECT 224.150 60.270 224.475 60.730 ;
        RECT 224.645 60.440 225.030 61.410 ;
        RECT 225.200 62.080 225.640 62.640 ;
        RECT 225.810 62.080 226.260 62.820 ;
        RECT 226.430 62.250 226.600 62.650 ;
        RECT 226.770 62.420 227.190 62.820 ;
        RECT 227.360 62.250 227.590 62.650 ;
        RECT 226.430 62.080 227.590 62.250 ;
        RECT 227.760 62.080 228.250 62.650 ;
        RECT 225.200 61.070 225.510 62.080 ;
        RECT 225.680 61.460 225.850 61.910 ;
        RECT 226.020 61.630 226.410 61.910 ;
        RECT 226.595 61.580 226.840 61.910 ;
        RECT 225.680 61.290 226.470 61.460 ;
        RECT 225.200 60.440 225.640 61.070 ;
        RECT 225.815 60.270 226.130 61.120 ;
        RECT 226.300 60.610 226.470 61.290 ;
        RECT 226.640 60.780 226.840 61.580 ;
        RECT 227.040 60.780 227.290 61.910 ;
        RECT 227.505 61.580 227.910 61.910 ;
        RECT 228.080 61.410 228.250 62.080 ;
        RECT 227.480 61.240 228.250 61.410 ;
        RECT 228.885 62.080 229.140 62.650 ;
        RECT 229.310 62.420 229.640 62.820 ;
        RECT 230.065 62.285 230.595 62.650 ;
        RECT 230.065 62.250 230.240 62.285 ;
        RECT 229.310 62.080 230.240 62.250 ;
        RECT 228.885 61.410 229.055 62.080 ;
        RECT 229.310 61.910 229.480 62.080 ;
        RECT 229.225 61.580 229.480 61.910 ;
        RECT 229.705 61.580 229.900 61.910 ;
        RECT 227.480 60.610 227.730 61.240 ;
        RECT 226.300 60.440 227.730 60.610 ;
        RECT 227.910 60.270 228.240 61.070 ;
        RECT 228.885 60.440 229.220 61.410 ;
        RECT 229.390 60.270 229.560 61.410 ;
        RECT 229.730 60.610 229.900 61.580 ;
        RECT 230.070 60.950 230.240 62.080 ;
        RECT 230.410 61.290 230.580 62.090 ;
        RECT 230.785 61.800 231.060 62.650 ;
        RECT 230.780 61.630 231.060 61.800 ;
        RECT 230.785 61.490 231.060 61.630 ;
        RECT 231.230 61.290 231.420 62.650 ;
        RECT 231.600 62.285 232.110 62.820 ;
        RECT 232.330 62.010 232.575 62.615 ;
        RECT 233.025 62.080 233.280 62.650 ;
        RECT 233.450 62.420 233.780 62.820 ;
        RECT 234.205 62.285 234.735 62.650 ;
        RECT 234.925 62.480 235.200 62.650 ;
        RECT 234.920 62.310 235.200 62.480 ;
        RECT 234.205 62.250 234.380 62.285 ;
        RECT 233.450 62.080 234.380 62.250 ;
        RECT 231.620 61.840 232.850 62.010 ;
        RECT 230.410 61.120 231.420 61.290 ;
        RECT 231.590 61.275 232.340 61.465 ;
        RECT 230.070 60.780 231.195 60.950 ;
        RECT 231.590 60.610 231.760 61.275 ;
        RECT 232.510 61.030 232.850 61.840 ;
        RECT 229.730 60.440 231.760 60.610 ;
        RECT 231.930 60.270 232.100 61.030 ;
        RECT 232.335 60.620 232.850 61.030 ;
        RECT 233.025 61.410 233.195 62.080 ;
        RECT 233.450 61.910 233.620 62.080 ;
        RECT 233.365 61.580 233.620 61.910 ;
        RECT 233.845 61.580 234.040 61.910 ;
        RECT 233.025 60.440 233.360 61.410 ;
        RECT 233.530 60.270 233.700 61.410 ;
        RECT 233.870 60.610 234.040 61.580 ;
        RECT 234.210 60.950 234.380 62.080 ;
        RECT 234.550 61.290 234.720 62.090 ;
        RECT 234.925 61.490 235.200 62.310 ;
        RECT 235.370 61.290 235.560 62.650 ;
        RECT 235.740 62.285 236.250 62.820 ;
        RECT 236.470 62.010 236.715 62.615 ;
        RECT 237.160 62.050 238.830 62.820 ;
        RECT 239.460 62.095 239.750 62.820 ;
        RECT 240.005 62.250 240.180 62.650 ;
        RECT 240.350 62.440 240.680 62.820 ;
        RECT 240.925 62.320 241.155 62.650 ;
        RECT 240.005 62.080 240.635 62.250 ;
        RECT 235.760 61.840 236.990 62.010 ;
        RECT 234.550 61.120 235.560 61.290 ;
        RECT 235.730 61.275 236.480 61.465 ;
        RECT 234.210 60.780 235.335 60.950 ;
        RECT 235.730 60.610 235.900 61.275 ;
        RECT 236.650 61.030 236.990 61.840 ;
        RECT 237.160 61.530 237.910 62.050 ;
        RECT 240.465 61.910 240.635 62.080 ;
        RECT 238.080 61.360 238.830 61.880 ;
        RECT 233.870 60.440 235.900 60.610 ;
        RECT 236.070 60.270 236.240 61.030 ;
        RECT 236.475 60.620 236.990 61.030 ;
        RECT 237.160 60.270 238.830 61.360 ;
        RECT 239.460 60.270 239.750 61.435 ;
        RECT 239.920 61.230 240.285 61.910 ;
        RECT 240.465 61.580 240.815 61.910 ;
        RECT 240.465 61.060 240.635 61.580 ;
        RECT 240.005 60.890 240.635 61.060 ;
        RECT 240.985 61.030 241.155 62.320 ;
        RECT 241.355 61.210 241.635 62.485 ;
        RECT 241.860 62.480 242.130 62.485 ;
        RECT 241.820 62.310 242.130 62.480 ;
        RECT 242.590 62.440 242.920 62.820 ;
        RECT 243.090 62.565 243.425 62.610 ;
        RECT 241.860 61.210 242.130 62.310 ;
        RECT 242.320 61.210 242.660 62.240 ;
        RECT 243.090 62.100 243.430 62.565 ;
        RECT 242.830 61.580 243.090 61.910 ;
        RECT 242.830 61.030 243.000 61.580 ;
        RECT 243.260 61.410 243.430 62.100 ;
        RECT 240.005 60.440 240.180 60.890 ;
        RECT 240.985 60.860 243.000 61.030 ;
        RECT 240.350 60.270 240.680 60.710 ;
        RECT 240.985 60.440 241.155 60.860 ;
        RECT 241.390 60.270 242.060 60.680 ;
        RECT 242.275 60.440 242.445 60.860 ;
        RECT 242.645 60.270 242.975 60.680 ;
        RECT 243.170 60.440 243.430 61.410 ;
        RECT 243.600 62.320 243.860 62.650 ;
        RECT 244.070 62.340 244.345 62.820 ;
        RECT 243.600 61.410 243.770 62.320 ;
        RECT 244.555 62.250 244.760 62.650 ;
        RECT 244.930 62.420 245.265 62.820 ;
        RECT 245.530 62.270 245.700 62.650 ;
        RECT 245.880 62.440 246.210 62.820 ;
        RECT 243.940 61.580 244.300 62.160 ;
        RECT 244.555 62.080 245.240 62.250 ;
        RECT 245.530 62.100 246.195 62.270 ;
        RECT 246.390 62.145 246.650 62.650 ;
        RECT 244.480 61.410 244.730 61.910 ;
        RECT 243.600 61.240 244.730 61.410 ;
        RECT 243.600 60.470 243.870 61.240 ;
        RECT 244.900 61.050 245.240 62.080 ;
        RECT 245.460 61.550 245.800 61.920 ;
        RECT 246.025 61.845 246.195 62.100 ;
        RECT 246.025 61.515 246.300 61.845 ;
        RECT 246.025 61.370 246.195 61.515 ;
        RECT 244.040 60.270 244.370 61.050 ;
        RECT 244.575 60.875 245.240 61.050 ;
        RECT 245.520 61.200 246.195 61.370 ;
        RECT 246.470 61.345 246.650 62.145 ;
        RECT 246.910 62.270 247.080 62.650 ;
        RECT 247.260 62.440 247.590 62.820 ;
        RECT 246.910 62.100 247.575 62.270 ;
        RECT 247.770 62.145 248.030 62.650 ;
        RECT 246.840 61.550 247.180 61.920 ;
        RECT 247.405 61.845 247.575 62.100 ;
        RECT 247.405 61.515 247.680 61.845 ;
        RECT 247.405 61.370 247.575 61.515 ;
        RECT 244.575 60.470 244.760 60.875 ;
        RECT 244.930 60.270 245.265 60.695 ;
        RECT 245.520 60.440 245.700 61.200 ;
        RECT 245.880 60.270 246.210 61.030 ;
        RECT 246.380 60.440 246.650 61.345 ;
        RECT 246.900 61.200 247.575 61.370 ;
        RECT 247.850 61.345 248.030 62.145 ;
        RECT 248.200 62.050 250.790 62.820 ;
        RECT 248.200 61.530 249.410 62.050 ;
        RECT 251.235 62.010 251.480 62.615 ;
        RECT 251.700 62.285 252.210 62.820 ;
        RECT 249.580 61.360 250.790 61.880 ;
        RECT 246.900 60.440 247.080 61.200 ;
        RECT 247.260 60.270 247.590 61.030 ;
        RECT 247.760 60.440 248.030 61.345 ;
        RECT 248.200 60.270 250.790 61.360 ;
        RECT 250.960 61.840 252.190 62.010 ;
        RECT 250.960 61.030 251.300 61.840 ;
        RECT 251.470 61.275 252.220 61.465 ;
        RECT 250.960 60.620 251.475 61.030 ;
        RECT 251.710 60.270 251.880 61.030 ;
        RECT 252.050 60.610 252.220 61.275 ;
        RECT 252.390 61.290 252.580 62.650 ;
        RECT 252.750 61.800 253.025 62.650 ;
        RECT 253.215 62.285 253.745 62.650 ;
        RECT 254.170 62.420 254.500 62.820 ;
        RECT 253.570 62.250 253.745 62.285 ;
        RECT 252.750 61.630 253.030 61.800 ;
        RECT 252.750 61.490 253.025 61.630 ;
        RECT 253.230 61.290 253.400 62.090 ;
        RECT 252.390 61.120 253.400 61.290 ;
        RECT 253.570 62.080 254.500 62.250 ;
        RECT 254.670 62.080 254.925 62.650 ;
        RECT 253.570 60.950 253.740 62.080 ;
        RECT 254.330 61.910 254.500 62.080 ;
        RECT 252.615 60.780 253.740 60.950 ;
        RECT 253.910 61.580 254.105 61.910 ;
        RECT 254.330 61.580 254.585 61.910 ;
        RECT 253.910 60.610 254.080 61.580 ;
        RECT 254.755 61.410 254.925 62.080 ;
        RECT 252.050 60.440 254.080 60.610 ;
        RECT 254.250 60.270 254.420 61.410 ;
        RECT 254.590 60.440 254.925 61.410 ;
        RECT 255.105 62.080 255.360 62.650 ;
        RECT 255.530 62.420 255.860 62.820 ;
        RECT 256.285 62.285 256.815 62.650 ;
        RECT 257.005 62.480 257.280 62.650 ;
        RECT 257.000 62.310 257.280 62.480 ;
        RECT 256.285 62.250 256.460 62.285 ;
        RECT 255.530 62.080 256.460 62.250 ;
        RECT 255.105 61.410 255.275 62.080 ;
        RECT 255.530 61.910 255.700 62.080 ;
        RECT 255.445 61.580 255.700 61.910 ;
        RECT 255.925 61.580 256.120 61.910 ;
        RECT 255.105 60.440 255.440 61.410 ;
        RECT 255.610 60.270 255.780 61.410 ;
        RECT 255.950 60.610 256.120 61.580 ;
        RECT 256.290 60.950 256.460 62.080 ;
        RECT 256.630 61.290 256.800 62.090 ;
        RECT 257.005 61.490 257.280 62.310 ;
        RECT 257.450 61.290 257.640 62.650 ;
        RECT 257.820 62.285 258.330 62.820 ;
        RECT 258.550 62.010 258.795 62.615 ;
        RECT 259.240 62.160 259.505 62.820 ;
        RECT 259.675 62.190 259.920 62.650 ;
        RECT 260.095 62.325 260.425 62.820 ;
        RECT 257.840 61.840 259.070 62.010 ;
        RECT 259.675 61.980 259.845 62.190 ;
        RECT 260.615 62.140 260.825 62.600 ;
        RECT 256.630 61.120 257.640 61.290 ;
        RECT 257.810 61.275 258.560 61.465 ;
        RECT 256.290 60.780 257.415 60.950 ;
        RECT 257.810 60.610 257.980 61.275 ;
        RECT 258.730 61.030 259.070 61.840 ;
        RECT 259.240 61.460 259.845 61.980 ;
        RECT 255.950 60.440 257.980 60.610 ;
        RECT 258.150 60.270 258.320 61.030 ;
        RECT 258.555 60.620 259.070 61.030 ;
        RECT 259.240 60.270 259.505 61.280 ;
        RECT 259.675 61.110 259.845 61.460 ;
        RECT 260.015 61.480 260.245 61.910 ;
        RECT 260.415 61.660 260.825 62.140 ;
        RECT 260.995 62.335 261.780 62.600 ;
        RECT 260.995 61.480 261.250 62.335 ;
        RECT 261.980 61.890 262.255 62.600 ;
        RECT 262.480 62.330 262.750 62.820 ;
        RECT 261.420 61.660 262.255 61.890 ;
        RECT 260.015 61.310 261.785 61.480 ;
        RECT 259.675 60.440 259.960 61.110 ;
        RECT 260.160 60.270 260.375 61.115 ;
        RECT 260.635 61.015 260.825 61.310 ;
        RECT 261.050 60.950 261.380 61.140 ;
        RECT 260.545 60.440 261.020 60.780 ;
        RECT 261.190 60.775 261.380 60.950 ;
        RECT 261.550 60.945 261.785 61.310 ;
        RECT 261.980 61.000 262.255 61.660 ;
        RECT 262.425 61.580 262.690 62.160 ;
        RECT 262.920 62.050 264.590 62.820 ;
        RECT 265.220 62.095 265.510 62.820 ;
        RECT 265.680 62.275 271.025 62.820 ;
        RECT 271.200 62.275 276.545 62.820 ;
        RECT 262.920 61.530 263.670 62.050 ;
        RECT 263.840 61.360 264.590 61.880 ;
        RECT 267.265 61.445 267.605 62.275 ;
        RECT 261.190 60.270 261.805 60.775 ;
        RECT 262.435 60.270 262.750 61.330 ;
        RECT 262.920 60.270 264.590 61.360 ;
        RECT 265.220 60.270 265.510 61.435 ;
        RECT 269.085 60.705 269.435 61.955 ;
        RECT 272.785 61.445 273.125 62.275 ;
        RECT 276.720 62.050 279.310 62.820 ;
        RECT 279.480 62.190 279.820 62.650 ;
        RECT 279.990 62.360 280.160 62.820 ;
        RECT 280.790 62.385 281.150 62.650 ;
        RECT 280.795 62.380 281.150 62.385 ;
        RECT 280.800 62.370 281.150 62.380 ;
        RECT 280.805 62.365 281.150 62.370 ;
        RECT 280.810 62.355 281.150 62.365 ;
        RECT 281.390 62.360 281.560 62.820 ;
        RECT 280.815 62.350 281.150 62.355 ;
        RECT 280.825 62.340 281.150 62.350 ;
        RECT 280.835 62.330 281.150 62.340 ;
        RECT 280.330 62.190 280.660 62.270 ;
        RECT 274.605 60.705 274.955 61.955 ;
        RECT 276.720 61.530 277.930 62.050 ;
        RECT 279.480 62.000 280.660 62.190 ;
        RECT 280.850 62.190 281.150 62.330 ;
        RECT 280.850 62.000 281.560 62.190 ;
        RECT 278.100 61.360 279.310 61.880 ;
        RECT 265.680 60.270 271.025 60.705 ;
        RECT 271.200 60.270 276.545 60.705 ;
        RECT 276.720 60.270 279.310 61.360 ;
        RECT 279.480 61.630 279.810 61.830 ;
        RECT 280.120 61.810 280.450 61.830 ;
        RECT 280.000 61.630 280.450 61.810 ;
        RECT 279.480 61.290 279.710 61.630 ;
        RECT 279.490 60.270 279.820 60.990 ;
        RECT 280.000 60.515 280.215 61.630 ;
        RECT 280.620 61.600 281.090 61.830 ;
        RECT 281.275 61.430 281.560 62.000 ;
        RECT 281.730 61.875 282.070 62.650 ;
        RECT 280.410 61.215 281.560 61.430 ;
        RECT 280.410 60.440 280.740 61.215 ;
        RECT 280.910 60.270 281.620 61.045 ;
        RECT 281.790 60.440 282.070 61.875 ;
        RECT 282.245 62.080 282.500 62.650 ;
        RECT 282.670 62.420 283.000 62.820 ;
        RECT 283.425 62.285 283.955 62.650 ;
        RECT 284.145 62.480 284.420 62.650 ;
        RECT 284.140 62.310 284.420 62.480 ;
        RECT 283.425 62.250 283.600 62.285 ;
        RECT 282.670 62.080 283.600 62.250 ;
        RECT 282.245 61.410 282.415 62.080 ;
        RECT 282.670 61.910 282.840 62.080 ;
        RECT 282.585 61.580 282.840 61.910 ;
        RECT 283.065 61.580 283.260 61.910 ;
        RECT 282.245 60.440 282.580 61.410 ;
        RECT 282.750 60.270 282.920 61.410 ;
        RECT 283.090 60.610 283.260 61.580 ;
        RECT 283.430 60.950 283.600 62.080 ;
        RECT 283.770 61.290 283.940 62.090 ;
        RECT 284.145 61.490 284.420 62.310 ;
        RECT 284.590 61.290 284.780 62.650 ;
        RECT 284.960 62.285 285.470 62.820 ;
        RECT 285.690 62.010 285.935 62.615 ;
        RECT 286.385 62.080 286.640 62.650 ;
        RECT 286.810 62.420 287.140 62.820 ;
        RECT 287.565 62.285 288.095 62.650 ;
        RECT 287.565 62.250 287.740 62.285 ;
        RECT 286.810 62.080 287.740 62.250 ;
        RECT 284.980 61.840 286.210 62.010 ;
        RECT 283.770 61.120 284.780 61.290 ;
        RECT 284.950 61.275 285.700 61.465 ;
        RECT 283.430 60.780 284.555 60.950 ;
        RECT 284.950 60.610 285.120 61.275 ;
        RECT 285.870 61.030 286.210 61.840 ;
        RECT 283.090 60.440 285.120 60.610 ;
        RECT 285.290 60.270 285.460 61.030 ;
        RECT 285.695 60.620 286.210 61.030 ;
        RECT 286.385 61.410 286.555 62.080 ;
        RECT 286.810 61.910 286.980 62.080 ;
        RECT 286.725 61.580 286.980 61.910 ;
        RECT 287.205 61.580 287.400 61.910 ;
        RECT 286.385 60.440 286.720 61.410 ;
        RECT 286.890 60.270 287.060 61.410 ;
        RECT 287.230 60.610 287.400 61.580 ;
        RECT 287.570 60.950 287.740 62.080 ;
        RECT 287.910 61.290 288.080 62.090 ;
        RECT 288.285 61.800 288.560 62.650 ;
        RECT 288.280 61.630 288.560 61.800 ;
        RECT 288.285 61.490 288.560 61.630 ;
        RECT 288.730 61.290 288.920 62.650 ;
        RECT 289.100 62.285 289.610 62.820 ;
        RECT 289.830 62.010 290.075 62.615 ;
        RECT 290.980 62.095 291.270 62.820 ;
        RECT 291.440 62.050 294.950 62.820 ;
        RECT 295.125 62.080 295.380 62.650 ;
        RECT 295.550 62.420 295.880 62.820 ;
        RECT 296.305 62.285 296.835 62.650 ;
        RECT 296.305 62.250 296.480 62.285 ;
        RECT 295.550 62.080 296.480 62.250 ;
        RECT 297.025 62.140 297.300 62.650 ;
        RECT 289.120 61.840 290.350 62.010 ;
        RECT 287.910 61.120 288.920 61.290 ;
        RECT 289.090 61.275 289.840 61.465 ;
        RECT 287.570 60.780 288.695 60.950 ;
        RECT 289.090 60.610 289.260 61.275 ;
        RECT 290.010 61.030 290.350 61.840 ;
        RECT 291.440 61.530 293.090 62.050 ;
        RECT 287.230 60.440 289.260 60.610 ;
        RECT 289.430 60.270 289.600 61.030 ;
        RECT 289.835 60.620 290.350 61.030 ;
        RECT 290.980 60.270 291.270 61.435 ;
        RECT 293.260 61.360 294.950 61.880 ;
        RECT 291.440 60.270 294.950 61.360 ;
        RECT 295.125 61.410 295.295 62.080 ;
        RECT 295.550 61.910 295.720 62.080 ;
        RECT 295.465 61.580 295.720 61.910 ;
        RECT 295.945 61.580 296.140 61.910 ;
        RECT 295.125 60.440 295.460 61.410 ;
        RECT 295.630 60.270 295.800 61.410 ;
        RECT 295.970 60.610 296.140 61.580 ;
        RECT 296.310 60.950 296.480 62.080 ;
        RECT 296.650 61.290 296.820 62.090 ;
        RECT 297.020 61.970 297.300 62.140 ;
        RECT 297.025 61.490 297.300 61.970 ;
        RECT 297.470 61.290 297.660 62.650 ;
        RECT 297.840 62.285 298.350 62.820 ;
        RECT 298.570 62.010 298.815 62.615 ;
        RECT 299.265 62.080 299.520 62.650 ;
        RECT 299.690 62.420 300.020 62.820 ;
        RECT 300.445 62.285 300.975 62.650 ;
        RECT 300.445 62.250 300.620 62.285 ;
        RECT 299.690 62.080 300.620 62.250 ;
        RECT 297.860 61.840 299.090 62.010 ;
        RECT 296.650 61.120 297.660 61.290 ;
        RECT 297.830 61.275 298.580 61.465 ;
        RECT 296.310 60.780 297.435 60.950 ;
        RECT 297.830 60.610 298.000 61.275 ;
        RECT 298.750 61.030 299.090 61.840 ;
        RECT 295.970 60.440 298.000 60.610 ;
        RECT 298.170 60.270 298.340 61.030 ;
        RECT 298.575 60.620 299.090 61.030 ;
        RECT 299.265 61.410 299.435 62.080 ;
        RECT 299.690 61.910 299.860 62.080 ;
        RECT 299.605 61.580 299.860 61.910 ;
        RECT 300.085 61.580 300.280 61.910 ;
        RECT 299.265 60.440 299.600 61.410 ;
        RECT 299.770 60.270 299.940 61.410 ;
        RECT 300.110 60.610 300.280 61.580 ;
        RECT 300.450 60.950 300.620 62.080 ;
        RECT 300.790 61.290 300.960 62.090 ;
        RECT 301.165 61.800 301.440 62.650 ;
        RECT 301.160 61.630 301.440 61.800 ;
        RECT 301.165 61.490 301.440 61.630 ;
        RECT 301.610 61.290 301.800 62.650 ;
        RECT 301.980 62.285 302.490 62.820 ;
        RECT 302.710 62.010 302.955 62.615 ;
        RECT 303.460 62.340 303.740 62.820 ;
        RECT 303.910 62.170 304.170 62.560 ;
        RECT 304.345 62.340 304.600 62.820 ;
        RECT 304.770 62.170 305.065 62.560 ;
        RECT 305.245 62.340 305.520 62.820 ;
        RECT 305.690 62.320 305.990 62.650 ;
        RECT 302.000 61.840 303.230 62.010 ;
        RECT 300.790 61.120 301.800 61.290 ;
        RECT 301.970 61.275 302.720 61.465 ;
        RECT 300.450 60.780 301.575 60.950 ;
        RECT 301.970 60.610 302.140 61.275 ;
        RECT 302.890 61.030 303.230 61.840 ;
        RECT 303.415 62.000 305.065 62.170 ;
        RECT 303.415 61.490 303.820 62.000 ;
        RECT 303.990 61.660 305.130 61.830 ;
        RECT 303.415 61.320 304.170 61.490 ;
        RECT 300.110 60.440 302.140 60.610 ;
        RECT 302.310 60.270 302.480 61.030 ;
        RECT 302.715 60.620 303.230 61.030 ;
        RECT 303.455 60.270 303.740 61.140 ;
        RECT 303.910 61.070 304.170 61.320 ;
        RECT 304.960 61.410 305.130 61.660 ;
        RECT 305.300 61.580 305.650 62.150 ;
        RECT 305.820 61.410 305.990 62.320 ;
        RECT 306.160 62.050 309.670 62.820 ;
        RECT 309.840 62.070 311.050 62.820 ;
        RECT 306.160 61.530 307.810 62.050 ;
        RECT 304.960 61.240 305.990 61.410 ;
        RECT 307.980 61.360 309.670 61.880 ;
        RECT 303.910 60.900 305.030 61.070 ;
        RECT 303.910 60.440 304.170 60.900 ;
        RECT 304.345 60.270 304.600 60.730 ;
        RECT 304.770 60.440 305.030 60.900 ;
        RECT 305.200 60.270 305.510 61.070 ;
        RECT 305.680 60.440 305.990 61.240 ;
        RECT 306.160 60.270 309.670 61.360 ;
        RECT 309.840 61.360 310.360 61.900 ;
        RECT 310.530 61.530 311.050 62.070 ;
        RECT 309.840 60.270 311.050 61.360 ;
        RECT 162.095 60.100 311.135 60.270 ;
        RECT 162.180 59.010 163.390 60.100 ;
        RECT 163.560 59.665 168.905 60.100 ;
        RECT 169.080 59.665 174.425 60.100 ;
        RECT 162.180 58.300 162.700 58.840 ;
        RECT 162.870 58.470 163.390 59.010 ;
        RECT 162.180 57.550 163.390 58.300 ;
        RECT 165.145 58.095 165.485 58.925 ;
        RECT 166.965 58.415 167.315 59.665 ;
        RECT 170.665 58.095 171.005 58.925 ;
        RECT 172.485 58.415 172.835 59.665 ;
        RECT 175.060 58.935 175.350 60.100 ;
        RECT 176.440 58.960 176.730 60.100 ;
        RECT 176.900 59.380 177.350 59.930 ;
        RECT 177.540 59.380 177.870 60.100 ;
        RECT 163.560 57.550 168.905 58.095 ;
        RECT 169.080 57.550 174.425 58.095 ;
        RECT 175.060 57.550 175.350 58.275 ;
        RECT 176.440 57.550 176.730 58.350 ;
        RECT 176.900 58.010 177.150 59.380 ;
        RECT 178.080 59.210 178.380 59.760 ;
        RECT 178.550 59.430 178.830 60.100 ;
        RECT 177.440 59.040 178.380 59.210 ;
        RECT 177.440 58.790 177.610 59.040 ;
        RECT 178.715 58.790 179.030 59.230 ;
        RECT 179.200 59.010 180.870 60.100 ;
        RECT 181.500 59.505 181.760 59.685 ;
        RECT 181.965 59.675 182.325 60.100 ;
        RECT 182.835 59.675 183.165 60.100 ;
        RECT 183.670 59.675 184.010 60.100 ;
        RECT 184.935 59.675 185.470 59.890 ;
        RECT 181.500 59.335 185.035 59.505 ;
        RECT 181.500 59.275 182.180 59.335 ;
        RECT 177.320 58.460 177.610 58.790 ;
        RECT 177.780 58.540 178.110 58.790 ;
        RECT 178.340 58.540 179.030 58.790 ;
        RECT 177.440 58.370 177.610 58.460 ;
        RECT 177.440 58.180 178.830 58.370 ;
        RECT 176.900 57.720 177.450 58.010 ;
        RECT 177.620 57.550 177.870 58.010 ;
        RECT 178.500 57.820 178.830 58.180 ;
        RECT 179.200 58.320 179.950 58.840 ;
        RECT 180.120 58.490 180.870 59.010 ;
        RECT 181.500 58.540 181.840 59.105 ;
        RECT 182.010 58.370 182.180 59.275 ;
        RECT 179.200 57.550 180.870 58.320 ;
        RECT 181.500 58.200 182.180 58.370 ;
        RECT 182.350 58.880 183.635 59.165 ;
        RECT 183.815 58.880 184.135 59.165 ;
        RECT 182.350 58.370 182.520 58.880 ;
        RECT 182.690 58.540 183.780 58.710 ;
        RECT 182.350 58.200 183.440 58.370 ;
        RECT 181.500 57.755 181.760 58.200 ;
        RECT 182.035 57.550 182.205 58.030 ;
        RECT 182.415 57.750 182.745 58.200 ;
        RECT 183.270 58.050 183.440 58.200 ;
        RECT 183.610 58.355 183.780 58.540 ;
        RECT 183.950 58.460 184.135 58.880 ;
        RECT 184.305 58.460 184.615 59.165 ;
        RECT 184.805 58.790 185.035 59.335 ;
        RECT 184.805 58.460 185.095 58.790 ;
        RECT 183.610 58.290 183.815 58.355 ;
        RECT 185.265 58.290 185.470 59.675 ;
        RECT 185.640 59.400 186.000 60.100 ;
        RECT 186.530 59.570 186.860 59.910 ;
        RECT 187.390 59.740 188.060 60.100 ;
        RECT 188.230 59.570 188.420 59.930 ;
        RECT 188.590 59.720 188.940 60.100 ;
        RECT 186.530 59.550 188.420 59.570 ;
        RECT 186.530 59.340 188.950 59.550 ;
        RECT 188.230 59.295 188.950 59.340 ;
        RECT 185.675 58.960 187.595 59.170 ;
        RECT 185.675 58.460 186.045 58.960 ;
        RECT 186.385 58.460 186.935 58.790 ;
        RECT 187.290 58.455 187.595 58.960 ;
        RECT 187.920 58.540 188.590 59.080 ;
        RECT 188.760 58.800 188.950 59.295 ;
        RECT 189.120 59.165 189.300 59.930 ;
        RECT 189.470 59.335 189.800 60.100 ;
        RECT 189.970 59.165 190.160 59.930 ;
        RECT 190.330 59.335 190.660 60.100 ;
        RECT 191.160 59.760 192.340 59.930 ;
        RECT 189.120 58.995 190.985 59.165 ;
        RECT 188.760 58.460 190.585 58.800 ;
        RECT 188.760 58.335 188.960 58.460 ;
        RECT 183.610 58.185 185.470 58.290 ;
        RECT 183.665 58.120 185.470 58.185 ;
        RECT 182.915 57.550 183.085 58.030 ;
        RECT 183.270 57.720 183.505 58.050 ;
        RECT 183.675 57.550 184.005 57.950 ;
        RECT 184.175 57.770 184.345 58.120 ;
        RECT 185.075 58.070 185.470 58.120 ;
        RECT 185.670 58.080 187.800 58.250 ;
        RECT 187.980 58.120 188.960 58.335 ;
        RECT 190.755 58.270 190.985 58.995 ;
        RECT 191.160 58.960 191.500 59.760 ;
        RECT 191.670 58.790 191.905 59.515 ;
        RECT 192.075 59.130 192.340 59.760 ;
        RECT 192.510 59.300 193.210 60.100 ;
        RECT 192.075 58.960 193.165 59.130 ;
        RECT 191.160 58.540 191.500 58.790 ;
        RECT 191.670 58.540 192.130 58.790 ;
        RECT 192.300 58.540 192.775 58.790 ;
        RECT 192.945 58.710 193.165 58.960 ;
        RECT 193.420 59.090 193.670 59.930 ;
        RECT 193.840 59.260 194.090 60.100 ;
        RECT 194.260 59.090 194.510 59.930 ;
        RECT 194.680 59.260 194.930 60.100 ;
        RECT 195.500 59.430 195.780 60.100 ;
        RECT 193.420 58.920 195.130 59.090 ;
        RECT 193.980 58.910 194.150 58.920 ;
        RECT 192.945 58.540 194.670 58.710 ;
        RECT 192.945 58.370 193.165 58.540 ;
        RECT 194.840 58.370 195.130 58.920 ;
        RECT 195.300 58.790 195.615 59.230 ;
        RECT 195.950 59.210 196.250 59.760 ;
        RECT 196.460 59.380 196.790 60.100 ;
        RECT 196.980 59.380 197.430 59.930 ;
        RECT 195.950 59.040 196.890 59.210 ;
        RECT 196.720 58.790 196.890 59.040 ;
        RECT 195.300 58.540 195.990 58.790 ;
        RECT 196.220 58.540 196.550 58.790 ;
        RECT 196.720 58.460 197.010 58.790 ;
        RECT 196.720 58.370 196.890 58.460 ;
        RECT 189.360 58.100 190.985 58.270 ;
        RECT 191.160 58.190 193.165 58.370 ;
        RECT 193.380 58.200 195.130 58.370 ;
        RECT 189.360 58.080 190.480 58.100 ;
        RECT 184.515 57.550 184.905 57.950 ;
        RECT 185.075 57.770 185.330 58.070 ;
        RECT 187.470 57.950 187.800 58.080 ;
        RECT 186.100 57.550 186.430 57.910 ;
        RECT 186.960 57.550 187.300 57.910 ;
        RECT 187.470 57.720 188.740 57.950 ;
        RECT 188.930 57.550 189.260 57.930 ;
        RECT 189.790 57.550 190.120 57.910 ;
        RECT 190.650 57.550 190.980 57.930 ;
        RECT 191.160 57.720 191.500 58.190 ;
        RECT 191.670 57.550 191.840 58.020 ;
        RECT 192.010 57.720 192.340 58.190 ;
        RECT 192.510 57.550 193.210 58.020 ;
        RECT 193.380 57.730 193.710 58.200 ;
        RECT 193.880 57.550 194.050 58.020 ;
        RECT 194.220 57.730 194.550 58.200 ;
        RECT 195.500 58.180 196.890 58.370 ;
        RECT 194.720 57.550 194.890 58.020 ;
        RECT 195.500 57.820 195.830 58.180 ;
        RECT 197.180 58.010 197.430 59.380 ;
        RECT 197.600 58.960 197.890 60.100 ;
        RECT 198.060 59.010 200.650 60.100 ;
        RECT 196.460 57.550 196.710 58.010 ;
        RECT 196.880 57.720 197.430 58.010 ;
        RECT 197.600 57.550 197.890 58.350 ;
        RECT 198.060 58.320 199.270 58.840 ;
        RECT 199.440 58.490 200.650 59.010 ;
        RECT 200.820 58.935 201.110 60.100 ;
        RECT 201.280 59.300 201.720 59.930 ;
        RECT 198.060 57.550 200.650 58.320 ;
        RECT 201.280 58.290 201.590 59.300 ;
        RECT 201.895 59.250 202.210 60.100 ;
        RECT 202.380 59.760 203.810 59.930 ;
        RECT 202.380 59.080 202.550 59.760 ;
        RECT 201.760 58.910 202.550 59.080 ;
        RECT 201.760 58.460 201.930 58.910 ;
        RECT 202.720 58.790 202.920 59.590 ;
        RECT 202.100 58.460 202.490 58.740 ;
        RECT 202.675 58.460 202.920 58.790 ;
        RECT 203.120 58.460 203.370 59.590 ;
        RECT 203.560 59.130 203.810 59.760 ;
        RECT 203.990 59.300 204.320 60.100 ;
        RECT 204.500 59.665 209.845 60.100 ;
        RECT 203.560 58.960 204.330 59.130 ;
        RECT 203.585 58.460 203.990 58.790 ;
        RECT 204.160 58.290 204.330 58.960 ;
        RECT 200.820 57.550 201.110 58.275 ;
        RECT 201.280 57.730 201.720 58.290 ;
        RECT 201.890 57.550 202.340 58.290 ;
        RECT 202.510 58.120 203.670 58.290 ;
        RECT 202.510 57.720 202.680 58.120 ;
        RECT 202.850 57.550 203.270 57.950 ;
        RECT 203.440 57.720 203.670 58.120 ;
        RECT 203.840 57.720 204.330 58.290 ;
        RECT 206.085 58.095 206.425 58.925 ;
        RECT 207.905 58.415 208.255 59.665 ;
        RECT 210.020 59.010 212.610 60.100 ;
        RECT 212.785 59.430 213.040 59.930 ;
        RECT 213.210 59.600 213.540 60.100 ;
        RECT 212.785 59.260 213.535 59.430 ;
        RECT 210.020 58.320 211.230 58.840 ;
        RECT 211.400 58.490 212.610 59.010 ;
        RECT 212.785 58.440 213.135 59.090 ;
        RECT 204.500 57.550 209.845 58.095 ;
        RECT 210.020 57.550 212.610 58.320 ;
        RECT 213.305 58.270 213.535 59.260 ;
        RECT 212.785 58.100 213.535 58.270 ;
        RECT 212.785 57.810 213.040 58.100 ;
        RECT 213.210 57.550 213.540 57.930 ;
        RECT 213.710 57.810 213.880 59.930 ;
        RECT 214.050 59.130 214.375 59.915 ;
        RECT 214.545 59.640 214.795 60.100 ;
        RECT 214.965 59.600 215.215 59.930 ;
        RECT 215.430 59.600 216.110 59.930 ;
        RECT 214.965 59.470 215.135 59.600 ;
        RECT 214.740 59.300 215.135 59.470 ;
        RECT 214.110 58.080 214.570 59.130 ;
        RECT 214.740 57.940 214.910 59.300 ;
        RECT 215.305 59.040 215.770 59.430 ;
        RECT 215.080 58.230 215.430 58.850 ;
        RECT 215.600 58.450 215.770 59.040 ;
        RECT 215.940 58.820 216.110 59.600 ;
        RECT 216.280 59.500 216.450 59.840 ;
        RECT 216.685 59.670 217.015 60.100 ;
        RECT 217.185 59.500 217.355 59.840 ;
        RECT 217.650 59.640 218.020 60.100 ;
        RECT 216.280 59.330 217.355 59.500 ;
        RECT 218.190 59.470 218.360 59.930 ;
        RECT 218.595 59.590 219.465 59.930 ;
        RECT 219.635 59.640 219.885 60.100 ;
        RECT 217.800 59.300 218.360 59.470 ;
        RECT 217.800 59.160 217.970 59.300 ;
        RECT 216.470 58.990 217.970 59.160 ;
        RECT 218.665 59.130 219.125 59.420 ;
        RECT 215.940 58.650 217.630 58.820 ;
        RECT 215.600 58.230 215.955 58.450 ;
        RECT 216.125 57.940 216.295 58.650 ;
        RECT 216.500 58.230 217.290 58.480 ;
        RECT 217.460 58.470 217.630 58.650 ;
        RECT 217.800 58.300 217.970 58.990 ;
        RECT 214.240 57.550 214.570 57.910 ;
        RECT 214.740 57.770 215.235 57.940 ;
        RECT 215.440 57.770 216.295 57.940 ;
        RECT 217.170 57.550 217.500 58.010 ;
        RECT 217.710 57.910 217.970 58.300 ;
        RECT 218.160 59.120 219.125 59.130 ;
        RECT 219.295 59.210 219.465 59.590 ;
        RECT 220.055 59.550 220.225 59.840 ;
        RECT 220.405 59.720 220.735 60.100 ;
        RECT 220.055 59.380 220.855 59.550 ;
        RECT 218.160 58.960 218.835 59.120 ;
        RECT 219.295 59.040 220.515 59.210 ;
        RECT 218.160 58.170 218.370 58.960 ;
        RECT 219.295 58.950 219.465 59.040 ;
        RECT 218.540 58.170 218.890 58.790 ;
        RECT 219.060 58.780 219.465 58.950 ;
        RECT 219.060 58.000 219.230 58.780 ;
        RECT 219.400 58.330 219.620 58.610 ;
        RECT 219.800 58.500 220.340 58.870 ;
        RECT 220.685 58.790 220.855 59.380 ;
        RECT 221.075 58.960 221.380 60.100 ;
        RECT 221.550 58.910 221.805 59.790 ;
        RECT 220.685 58.760 221.425 58.790 ;
        RECT 219.400 58.160 219.930 58.330 ;
        RECT 217.710 57.740 218.060 57.910 ;
        RECT 218.280 57.720 219.230 58.000 ;
        RECT 219.400 57.550 219.590 57.990 ;
        RECT 219.760 57.930 219.930 58.160 ;
        RECT 220.100 58.100 220.340 58.500 ;
        RECT 220.510 58.460 221.425 58.760 ;
        RECT 220.510 58.285 220.835 58.460 ;
        RECT 220.510 57.930 220.830 58.285 ;
        RECT 221.595 58.260 221.805 58.910 ;
        RECT 219.760 57.760 220.830 57.930 ;
        RECT 221.075 57.550 221.380 58.010 ;
        RECT 221.550 57.730 221.805 58.260 ;
        RECT 221.985 58.960 222.320 59.930 ;
        RECT 222.490 58.960 222.660 60.100 ;
        RECT 222.830 59.760 224.860 59.930 ;
        RECT 221.985 58.290 222.155 58.960 ;
        RECT 222.830 58.790 223.000 59.760 ;
        RECT 222.325 58.460 222.580 58.790 ;
        RECT 222.805 58.460 223.000 58.790 ;
        RECT 223.170 59.420 224.295 59.590 ;
        RECT 222.410 58.290 222.580 58.460 ;
        RECT 223.170 58.290 223.340 59.420 ;
        RECT 221.985 57.720 222.240 58.290 ;
        RECT 222.410 58.120 223.340 58.290 ;
        RECT 223.510 59.080 224.520 59.250 ;
        RECT 223.510 58.280 223.680 59.080 ;
        RECT 223.885 58.400 224.160 58.880 ;
        RECT 223.880 58.230 224.160 58.400 ;
        RECT 223.165 58.085 223.340 58.120 ;
        RECT 222.410 57.550 222.740 57.950 ;
        RECT 223.165 57.720 223.695 58.085 ;
        RECT 223.885 57.720 224.160 58.230 ;
        RECT 224.330 57.720 224.520 59.080 ;
        RECT 224.690 59.095 224.860 59.760 ;
        RECT 225.030 59.340 225.200 60.100 ;
        RECT 225.435 59.340 225.950 59.750 ;
        RECT 224.690 58.905 225.440 59.095 ;
        RECT 225.610 58.530 225.950 59.340 ;
        RECT 226.580 58.935 226.870 60.100 ;
        RECT 227.615 59.470 227.900 59.930 ;
        RECT 228.070 59.640 228.340 60.100 ;
        RECT 227.615 59.250 228.570 59.470 ;
        RECT 224.720 58.360 225.950 58.530 ;
        RECT 227.500 58.520 228.190 59.080 ;
        RECT 224.700 57.550 225.210 58.085 ;
        RECT 225.430 57.755 225.675 58.360 ;
        RECT 228.360 58.350 228.570 59.250 ;
        RECT 226.580 57.550 226.870 58.275 ;
        RECT 227.615 58.180 228.570 58.350 ;
        RECT 228.740 59.080 229.140 59.930 ;
        RECT 229.330 59.470 229.610 59.930 ;
        RECT 230.130 59.640 230.455 60.100 ;
        RECT 229.330 59.250 230.455 59.470 ;
        RECT 228.740 58.520 229.835 59.080 ;
        RECT 230.005 58.790 230.455 59.250 ;
        RECT 230.625 58.960 231.010 59.930 ;
        RECT 231.185 59.430 231.440 59.930 ;
        RECT 231.610 59.600 231.940 60.100 ;
        RECT 231.185 59.260 231.935 59.430 ;
        RECT 227.615 57.720 227.900 58.180 ;
        RECT 228.070 57.550 228.340 58.010 ;
        RECT 228.740 57.720 229.140 58.520 ;
        RECT 230.005 58.460 230.560 58.790 ;
        RECT 230.005 58.350 230.455 58.460 ;
        RECT 229.330 58.180 230.455 58.350 ;
        RECT 230.730 58.290 231.010 58.960 ;
        RECT 231.185 58.440 231.535 59.090 ;
        RECT 229.330 57.720 229.610 58.180 ;
        RECT 230.130 57.550 230.455 58.010 ;
        RECT 230.625 57.720 231.010 58.290 ;
        RECT 231.705 58.270 231.935 59.260 ;
        RECT 231.185 58.100 231.935 58.270 ;
        RECT 231.185 57.810 231.440 58.100 ;
        RECT 231.610 57.550 231.940 57.930 ;
        RECT 232.110 57.810 232.280 59.930 ;
        RECT 232.450 59.130 232.775 59.915 ;
        RECT 232.945 59.640 233.195 60.100 ;
        RECT 233.365 59.600 233.615 59.930 ;
        RECT 233.830 59.600 234.510 59.930 ;
        RECT 233.365 59.470 233.535 59.600 ;
        RECT 233.140 59.300 233.535 59.470 ;
        RECT 232.510 58.080 232.970 59.130 ;
        RECT 233.140 57.940 233.310 59.300 ;
        RECT 233.705 59.040 234.170 59.430 ;
        RECT 233.480 58.230 233.830 58.850 ;
        RECT 234.000 58.450 234.170 59.040 ;
        RECT 234.340 58.820 234.510 59.600 ;
        RECT 234.680 59.500 234.850 59.840 ;
        RECT 235.085 59.670 235.415 60.100 ;
        RECT 235.585 59.500 235.755 59.840 ;
        RECT 236.050 59.640 236.420 60.100 ;
        RECT 234.680 59.330 235.755 59.500 ;
        RECT 236.590 59.470 236.760 59.930 ;
        RECT 236.995 59.590 237.865 59.930 ;
        RECT 238.035 59.640 238.285 60.100 ;
        RECT 236.200 59.300 236.760 59.470 ;
        RECT 236.200 59.160 236.370 59.300 ;
        RECT 234.870 58.990 236.370 59.160 ;
        RECT 237.065 59.130 237.525 59.420 ;
        RECT 234.340 58.650 236.030 58.820 ;
        RECT 234.000 58.230 234.355 58.450 ;
        RECT 234.525 57.940 234.695 58.650 ;
        RECT 234.900 58.230 235.690 58.480 ;
        RECT 235.860 58.470 236.030 58.650 ;
        RECT 236.200 58.300 236.370 58.990 ;
        RECT 232.640 57.550 232.970 57.910 ;
        RECT 233.140 57.770 233.635 57.940 ;
        RECT 233.840 57.770 234.695 57.940 ;
        RECT 235.570 57.550 235.900 58.010 ;
        RECT 236.110 57.910 236.370 58.300 ;
        RECT 236.560 59.120 237.525 59.130 ;
        RECT 237.695 59.210 237.865 59.590 ;
        RECT 238.455 59.550 238.625 59.840 ;
        RECT 238.805 59.720 239.135 60.100 ;
        RECT 238.455 59.380 239.255 59.550 ;
        RECT 236.560 58.960 237.235 59.120 ;
        RECT 237.695 59.040 238.915 59.210 ;
        RECT 236.560 58.170 236.770 58.960 ;
        RECT 237.695 58.950 237.865 59.040 ;
        RECT 236.940 58.170 237.290 58.790 ;
        RECT 237.460 58.780 237.865 58.950 ;
        RECT 237.460 58.000 237.630 58.780 ;
        RECT 237.800 58.330 238.020 58.610 ;
        RECT 238.200 58.500 238.740 58.870 ;
        RECT 239.085 58.790 239.255 59.380 ;
        RECT 239.475 58.960 239.780 60.100 ;
        RECT 239.950 58.910 240.205 59.790 ;
        RECT 240.380 59.010 242.050 60.100 ;
        RECT 242.305 59.480 242.480 59.930 ;
        RECT 242.650 59.660 242.980 60.100 ;
        RECT 243.285 59.510 243.455 59.930 ;
        RECT 243.690 59.690 244.360 60.100 ;
        RECT 244.575 59.510 244.745 59.930 ;
        RECT 244.945 59.690 245.275 60.100 ;
        RECT 242.305 59.310 242.935 59.480 ;
        RECT 239.085 58.760 239.825 58.790 ;
        RECT 237.800 58.160 238.330 58.330 ;
        RECT 236.110 57.740 236.460 57.910 ;
        RECT 236.680 57.720 237.630 58.000 ;
        RECT 237.800 57.550 237.990 57.990 ;
        RECT 238.160 57.930 238.330 58.160 ;
        RECT 238.500 58.100 238.740 58.500 ;
        RECT 238.910 58.460 239.825 58.760 ;
        RECT 238.910 58.285 239.235 58.460 ;
        RECT 238.910 57.930 239.230 58.285 ;
        RECT 239.995 58.260 240.205 58.910 ;
        RECT 238.160 57.760 239.230 57.930 ;
        RECT 239.475 57.550 239.780 58.010 ;
        RECT 239.950 57.730 240.205 58.260 ;
        RECT 240.380 58.320 241.130 58.840 ;
        RECT 241.300 58.490 242.050 59.010 ;
        RECT 242.220 58.460 242.585 59.140 ;
        RECT 242.765 58.790 242.935 59.310 ;
        RECT 243.285 59.340 245.300 59.510 ;
        RECT 242.765 58.460 243.115 58.790 ;
        RECT 240.380 57.550 242.050 58.320 ;
        RECT 242.765 58.290 242.935 58.460 ;
        RECT 242.305 58.120 242.935 58.290 ;
        RECT 242.305 57.720 242.480 58.120 ;
        RECT 243.285 58.050 243.455 59.340 ;
        RECT 242.650 57.550 242.980 57.930 ;
        RECT 243.225 57.720 243.455 58.050 ;
        RECT 243.655 57.885 243.935 59.160 ;
        RECT 244.160 58.060 244.430 59.160 ;
        RECT 244.620 58.130 244.960 59.160 ;
        RECT 245.130 58.790 245.300 59.340 ;
        RECT 245.470 58.960 245.730 59.930 ;
        RECT 245.900 59.665 251.245 60.100 ;
        RECT 245.130 58.460 245.390 58.790 ;
        RECT 245.560 58.270 245.730 58.960 ;
        RECT 244.120 57.890 244.430 58.060 ;
        RECT 244.160 57.885 244.430 57.890 ;
        RECT 244.890 57.550 245.220 57.930 ;
        RECT 245.390 57.805 245.730 58.270 ;
        RECT 247.485 58.095 247.825 58.925 ;
        RECT 249.305 58.415 249.655 59.665 ;
        RECT 252.340 58.935 252.630 60.100 ;
        RECT 252.805 59.430 253.060 59.930 ;
        RECT 253.230 59.600 253.560 60.100 ;
        RECT 252.805 59.260 253.555 59.430 ;
        RECT 252.805 58.440 253.155 59.090 ;
        RECT 245.390 57.760 245.725 57.805 ;
        RECT 245.900 57.550 251.245 58.095 ;
        RECT 252.340 57.550 252.630 58.275 ;
        RECT 253.325 58.270 253.555 59.260 ;
        RECT 252.805 58.100 253.555 58.270 ;
        RECT 252.805 57.810 253.060 58.100 ;
        RECT 253.230 57.550 253.560 57.930 ;
        RECT 253.730 57.810 253.900 59.930 ;
        RECT 254.070 59.130 254.395 59.915 ;
        RECT 254.565 59.640 254.815 60.100 ;
        RECT 254.985 59.600 255.235 59.930 ;
        RECT 255.450 59.600 256.130 59.930 ;
        RECT 254.985 59.470 255.155 59.600 ;
        RECT 254.760 59.300 255.155 59.470 ;
        RECT 254.130 58.080 254.590 59.130 ;
        RECT 254.760 57.940 254.930 59.300 ;
        RECT 255.325 59.040 255.790 59.430 ;
        RECT 255.100 58.230 255.450 58.850 ;
        RECT 255.620 58.450 255.790 59.040 ;
        RECT 255.960 58.820 256.130 59.600 ;
        RECT 256.300 59.500 256.470 59.840 ;
        RECT 256.705 59.670 257.035 60.100 ;
        RECT 257.205 59.500 257.375 59.840 ;
        RECT 257.670 59.640 258.040 60.100 ;
        RECT 256.300 59.330 257.375 59.500 ;
        RECT 258.210 59.470 258.380 59.930 ;
        RECT 258.615 59.590 259.485 59.930 ;
        RECT 259.655 59.640 259.905 60.100 ;
        RECT 257.820 59.300 258.380 59.470 ;
        RECT 257.820 59.160 257.990 59.300 ;
        RECT 256.490 58.990 257.990 59.160 ;
        RECT 258.685 59.130 259.145 59.420 ;
        RECT 255.960 58.650 257.650 58.820 ;
        RECT 255.620 58.230 255.975 58.450 ;
        RECT 256.145 57.940 256.315 58.650 ;
        RECT 256.520 58.230 257.310 58.480 ;
        RECT 257.480 58.470 257.650 58.650 ;
        RECT 257.820 58.300 257.990 58.990 ;
        RECT 254.260 57.550 254.590 57.910 ;
        RECT 254.760 57.770 255.255 57.940 ;
        RECT 255.460 57.770 256.315 57.940 ;
        RECT 257.190 57.550 257.520 58.010 ;
        RECT 257.730 57.910 257.990 58.300 ;
        RECT 258.180 59.120 259.145 59.130 ;
        RECT 259.315 59.210 259.485 59.590 ;
        RECT 260.075 59.550 260.245 59.840 ;
        RECT 260.425 59.720 260.755 60.100 ;
        RECT 260.075 59.380 260.875 59.550 ;
        RECT 258.180 58.960 258.855 59.120 ;
        RECT 259.315 59.040 260.535 59.210 ;
        RECT 258.180 58.170 258.390 58.960 ;
        RECT 259.315 58.950 259.485 59.040 ;
        RECT 258.560 58.170 258.910 58.790 ;
        RECT 259.080 58.780 259.485 58.950 ;
        RECT 259.080 58.000 259.250 58.780 ;
        RECT 259.420 58.330 259.640 58.610 ;
        RECT 259.820 58.500 260.360 58.870 ;
        RECT 260.705 58.790 260.875 59.380 ;
        RECT 261.095 58.960 261.400 60.100 ;
        RECT 261.570 58.910 261.825 59.790 ;
        RECT 260.705 58.760 261.445 58.790 ;
        RECT 259.420 58.160 259.950 58.330 ;
        RECT 257.730 57.740 258.080 57.910 ;
        RECT 258.300 57.720 259.250 58.000 ;
        RECT 259.420 57.550 259.610 57.990 ;
        RECT 259.780 57.930 259.950 58.160 ;
        RECT 260.120 58.100 260.360 58.500 ;
        RECT 260.530 58.460 261.445 58.760 ;
        RECT 260.530 58.285 260.855 58.460 ;
        RECT 260.530 57.930 260.850 58.285 ;
        RECT 261.615 58.260 261.825 58.910 ;
        RECT 259.780 57.760 260.850 57.930 ;
        RECT 261.095 57.550 261.400 58.010 ;
        RECT 261.570 57.730 261.825 58.260 ;
        RECT 262.000 59.670 262.340 59.930 ;
        RECT 262.000 58.270 262.260 59.670 ;
        RECT 262.510 59.300 262.840 60.100 ;
        RECT 263.305 59.130 263.555 59.930 ;
        RECT 263.740 59.380 264.070 60.100 ;
        RECT 264.290 59.130 264.540 59.930 ;
        RECT 264.710 59.720 265.045 60.100 ;
        RECT 262.450 58.960 264.640 59.130 ;
        RECT 262.450 58.790 262.765 58.960 ;
        RECT 262.435 58.540 262.765 58.790 ;
        RECT 262.000 57.760 262.340 58.270 ;
        RECT 262.510 57.550 262.780 58.350 ;
        RECT 262.960 57.820 263.240 58.790 ;
        RECT 263.420 57.820 263.720 58.790 ;
        RECT 263.900 57.825 264.250 58.790 ;
        RECT 264.470 58.050 264.640 58.960 ;
        RECT 264.810 58.230 265.050 59.540 ;
        RECT 265.220 59.010 268.730 60.100 ;
        RECT 268.900 59.010 270.110 60.100 ;
        RECT 270.960 59.740 271.290 60.100 ;
        RECT 271.815 59.740 272.150 60.100 ;
        RECT 272.720 59.740 273.050 60.100 ;
        RECT 273.615 59.740 274.065 60.100 ;
        RECT 265.220 58.320 266.870 58.840 ;
        RECT 267.040 58.490 268.730 59.010 ;
        RECT 264.470 57.720 264.965 58.050 ;
        RECT 265.220 57.550 268.730 58.320 ;
        RECT 268.900 58.300 269.420 58.840 ;
        RECT 269.590 58.470 270.110 59.010 ;
        RECT 270.350 59.340 274.115 59.570 ;
        RECT 268.900 57.550 270.110 58.300 ;
        RECT 270.350 57.890 270.630 59.340 ;
        RECT 270.800 58.080 271.080 59.170 ;
        RECT 271.260 59.000 272.570 59.170 ;
        RECT 271.260 58.310 271.525 59.000 ;
        RECT 272.740 58.990 273.515 59.160 ;
        RECT 272.740 58.820 272.910 58.990 ;
        RECT 271.695 58.485 272.910 58.820 ;
        RECT 271.260 58.080 272.510 58.310 ;
        RECT 272.680 58.270 272.910 58.485 ;
        RECT 273.080 58.460 273.270 58.805 ;
        RECT 272.680 58.080 273.375 58.270 ;
        RECT 273.560 58.190 273.775 58.805 ;
        RECT 273.945 58.790 274.115 59.340 ;
        RECT 274.285 58.960 274.645 59.630 ;
        RECT 274.880 59.010 277.470 60.100 ;
        RECT 273.945 58.460 274.255 58.790 ;
        RECT 274.425 58.270 274.645 58.960 ;
        RECT 270.960 57.550 271.290 57.910 ;
        RECT 271.460 57.720 271.650 58.080 ;
        RECT 272.320 57.980 272.510 58.080 ;
        RECT 273.195 58.010 273.375 58.080 ;
        RECT 274.160 58.010 274.645 58.270 ;
        RECT 271.820 57.550 272.150 57.910 ;
        RECT 272.685 57.550 273.015 57.910 ;
        RECT 273.195 57.820 274.645 58.010 ;
        RECT 274.160 57.720 274.645 57.820 ;
        RECT 274.880 58.320 276.090 58.840 ;
        RECT 276.260 58.490 277.470 59.010 ;
        RECT 278.100 58.935 278.390 60.100 ;
        RECT 278.565 58.960 278.900 59.930 ;
        RECT 279.070 58.960 279.240 60.100 ;
        RECT 279.410 59.760 281.440 59.930 ;
        RECT 274.880 57.550 277.470 58.320 ;
        RECT 278.565 58.290 278.735 58.960 ;
        RECT 279.410 58.790 279.580 59.760 ;
        RECT 278.905 58.460 279.160 58.790 ;
        RECT 279.385 58.460 279.580 58.790 ;
        RECT 279.750 59.420 280.875 59.590 ;
        RECT 278.990 58.290 279.160 58.460 ;
        RECT 279.750 58.290 279.920 59.420 ;
        RECT 278.100 57.550 278.390 58.275 ;
        RECT 278.565 57.720 278.820 58.290 ;
        RECT 278.990 58.120 279.920 58.290 ;
        RECT 280.090 59.080 281.100 59.250 ;
        RECT 280.090 58.280 280.260 59.080 ;
        RECT 280.465 58.740 280.740 58.880 ;
        RECT 280.460 58.570 280.740 58.740 ;
        RECT 279.745 58.085 279.920 58.120 ;
        RECT 278.990 57.550 279.320 57.950 ;
        RECT 279.745 57.720 280.275 58.085 ;
        RECT 280.465 57.720 280.740 58.570 ;
        RECT 280.910 57.720 281.100 59.080 ;
        RECT 281.270 59.095 281.440 59.760 ;
        RECT 281.610 59.340 281.780 60.100 ;
        RECT 282.015 59.340 282.530 59.750 ;
        RECT 281.270 58.905 282.020 59.095 ;
        RECT 282.190 58.530 282.530 59.340 ;
        RECT 283.165 59.430 283.420 59.930 ;
        RECT 283.590 59.600 283.920 60.100 ;
        RECT 283.165 59.260 283.915 59.430 ;
        RECT 281.300 58.360 282.530 58.530 ;
        RECT 283.165 58.440 283.515 59.090 ;
        RECT 281.280 57.550 281.790 58.085 ;
        RECT 282.010 57.755 282.255 58.360 ;
        RECT 283.685 58.270 283.915 59.260 ;
        RECT 283.165 58.100 283.915 58.270 ;
        RECT 283.165 57.810 283.420 58.100 ;
        RECT 283.590 57.550 283.920 57.930 ;
        RECT 284.090 57.810 284.260 59.930 ;
        RECT 284.430 59.130 284.755 59.915 ;
        RECT 284.925 59.640 285.175 60.100 ;
        RECT 285.345 59.600 285.595 59.930 ;
        RECT 285.810 59.600 286.490 59.930 ;
        RECT 285.345 59.470 285.515 59.600 ;
        RECT 285.120 59.300 285.515 59.470 ;
        RECT 284.490 58.080 284.950 59.130 ;
        RECT 285.120 57.940 285.290 59.300 ;
        RECT 285.685 59.040 286.150 59.430 ;
        RECT 285.460 58.230 285.810 58.850 ;
        RECT 285.980 58.450 286.150 59.040 ;
        RECT 286.320 58.820 286.490 59.600 ;
        RECT 286.660 59.500 286.830 59.840 ;
        RECT 287.065 59.670 287.395 60.100 ;
        RECT 287.565 59.500 287.735 59.840 ;
        RECT 288.030 59.640 288.400 60.100 ;
        RECT 286.660 59.330 287.735 59.500 ;
        RECT 288.570 59.470 288.740 59.930 ;
        RECT 288.975 59.590 289.845 59.930 ;
        RECT 290.015 59.640 290.265 60.100 ;
        RECT 288.180 59.300 288.740 59.470 ;
        RECT 288.180 59.160 288.350 59.300 ;
        RECT 286.850 58.990 288.350 59.160 ;
        RECT 289.045 59.130 289.505 59.420 ;
        RECT 286.320 58.650 288.010 58.820 ;
        RECT 285.980 58.230 286.335 58.450 ;
        RECT 286.505 57.940 286.675 58.650 ;
        RECT 286.880 58.230 287.670 58.480 ;
        RECT 287.840 58.470 288.010 58.650 ;
        RECT 288.180 58.300 288.350 58.990 ;
        RECT 284.620 57.550 284.950 57.910 ;
        RECT 285.120 57.770 285.615 57.940 ;
        RECT 285.820 57.770 286.675 57.940 ;
        RECT 287.550 57.550 287.880 58.010 ;
        RECT 288.090 57.910 288.350 58.300 ;
        RECT 288.540 59.120 289.505 59.130 ;
        RECT 289.675 59.210 289.845 59.590 ;
        RECT 290.435 59.550 290.605 59.840 ;
        RECT 290.785 59.720 291.115 60.100 ;
        RECT 290.435 59.380 291.235 59.550 ;
        RECT 288.540 58.960 289.215 59.120 ;
        RECT 289.675 59.040 290.895 59.210 ;
        RECT 288.540 58.170 288.750 58.960 ;
        RECT 289.675 58.950 289.845 59.040 ;
        RECT 288.920 58.170 289.270 58.790 ;
        RECT 289.440 58.780 289.845 58.950 ;
        RECT 289.440 58.000 289.610 58.780 ;
        RECT 289.780 58.330 290.000 58.610 ;
        RECT 290.180 58.500 290.720 58.870 ;
        RECT 291.065 58.790 291.235 59.380 ;
        RECT 291.455 58.960 291.760 60.100 ;
        RECT 291.930 58.910 292.180 59.790 ;
        RECT 292.350 58.960 292.600 60.100 ;
        RECT 292.820 59.010 294.490 60.100 ;
        RECT 291.065 58.760 291.805 58.790 ;
        RECT 289.780 58.160 290.310 58.330 ;
        RECT 288.090 57.740 288.440 57.910 ;
        RECT 288.660 57.720 289.610 58.000 ;
        RECT 289.780 57.550 289.970 57.990 ;
        RECT 290.140 57.930 290.310 58.160 ;
        RECT 290.480 58.100 290.720 58.500 ;
        RECT 290.890 58.460 291.805 58.760 ;
        RECT 290.890 58.285 291.215 58.460 ;
        RECT 290.890 57.930 291.210 58.285 ;
        RECT 291.975 58.260 292.180 58.910 ;
        RECT 292.820 58.320 293.570 58.840 ;
        RECT 293.740 58.490 294.490 59.010 ;
        RECT 294.665 58.910 294.920 59.790 ;
        RECT 295.090 58.960 295.395 60.100 ;
        RECT 295.735 59.720 296.065 60.100 ;
        RECT 296.245 59.550 296.415 59.840 ;
        RECT 296.585 59.640 296.835 60.100 ;
        RECT 295.615 59.380 296.415 59.550 ;
        RECT 297.005 59.590 297.875 59.930 ;
        RECT 290.140 57.760 291.210 57.930 ;
        RECT 291.455 57.550 291.760 58.010 ;
        RECT 291.930 57.730 292.180 58.260 ;
        RECT 292.350 57.550 292.600 58.305 ;
        RECT 292.820 57.550 294.490 58.320 ;
        RECT 294.665 58.260 294.875 58.910 ;
        RECT 295.615 58.790 295.785 59.380 ;
        RECT 297.005 59.210 297.175 59.590 ;
        RECT 298.110 59.470 298.280 59.930 ;
        RECT 298.450 59.640 298.820 60.100 ;
        RECT 299.115 59.500 299.285 59.840 ;
        RECT 299.455 59.670 299.785 60.100 ;
        RECT 300.020 59.500 300.190 59.840 ;
        RECT 295.955 59.040 297.175 59.210 ;
        RECT 297.345 59.130 297.805 59.420 ;
        RECT 298.110 59.300 298.670 59.470 ;
        RECT 299.115 59.330 300.190 59.500 ;
        RECT 300.360 59.600 301.040 59.930 ;
        RECT 301.255 59.600 301.505 59.930 ;
        RECT 301.675 59.640 301.925 60.100 ;
        RECT 298.500 59.160 298.670 59.300 ;
        RECT 297.345 59.120 298.310 59.130 ;
        RECT 297.005 58.950 297.175 59.040 ;
        RECT 297.635 58.960 298.310 59.120 ;
        RECT 295.045 58.760 295.785 58.790 ;
        RECT 295.045 58.460 295.960 58.760 ;
        RECT 295.635 58.285 295.960 58.460 ;
        RECT 294.665 57.730 294.920 58.260 ;
        RECT 295.090 57.550 295.395 58.010 ;
        RECT 295.640 57.930 295.960 58.285 ;
        RECT 296.130 58.500 296.670 58.870 ;
        RECT 297.005 58.780 297.410 58.950 ;
        RECT 296.130 58.100 296.370 58.500 ;
        RECT 296.850 58.330 297.070 58.610 ;
        RECT 296.540 58.160 297.070 58.330 ;
        RECT 296.540 57.930 296.710 58.160 ;
        RECT 297.240 58.000 297.410 58.780 ;
        RECT 297.580 58.170 297.930 58.790 ;
        RECT 298.100 58.170 298.310 58.960 ;
        RECT 298.500 58.990 300.000 59.160 ;
        RECT 298.500 58.300 298.670 58.990 ;
        RECT 300.360 58.820 300.530 59.600 ;
        RECT 301.335 59.470 301.505 59.600 ;
        RECT 298.840 58.650 300.530 58.820 ;
        RECT 300.700 59.040 301.165 59.430 ;
        RECT 301.335 59.300 301.730 59.470 ;
        RECT 298.840 58.470 299.010 58.650 ;
        RECT 295.640 57.760 296.710 57.930 ;
        RECT 296.880 57.550 297.070 57.990 ;
        RECT 297.240 57.720 298.190 58.000 ;
        RECT 298.500 57.910 298.760 58.300 ;
        RECT 299.180 58.230 299.970 58.480 ;
        RECT 298.410 57.740 298.760 57.910 ;
        RECT 298.970 57.550 299.300 58.010 ;
        RECT 300.175 57.940 300.345 58.650 ;
        RECT 300.700 58.450 300.870 59.040 ;
        RECT 300.515 58.230 300.870 58.450 ;
        RECT 301.040 58.230 301.390 58.850 ;
        RECT 301.560 57.940 301.730 59.300 ;
        RECT 302.095 59.130 302.420 59.915 ;
        RECT 301.900 58.080 302.360 59.130 ;
        RECT 300.175 57.770 301.030 57.940 ;
        RECT 301.235 57.770 301.730 57.940 ;
        RECT 301.900 57.550 302.230 57.910 ;
        RECT 302.590 57.810 302.760 59.930 ;
        RECT 302.930 59.600 303.260 60.100 ;
        RECT 303.430 59.430 303.685 59.930 ;
        RECT 302.935 59.260 303.685 59.430 ;
        RECT 302.935 58.270 303.165 59.260 ;
        RECT 303.335 58.440 303.685 59.090 ;
        RECT 303.860 58.935 304.150 60.100 ;
        RECT 304.320 59.665 309.665 60.100 ;
        RECT 302.935 58.100 303.685 58.270 ;
        RECT 302.930 57.550 303.260 57.930 ;
        RECT 303.430 57.810 303.685 58.100 ;
        RECT 303.860 57.550 304.150 58.275 ;
        RECT 305.905 58.095 306.245 58.925 ;
        RECT 307.725 58.415 308.075 59.665 ;
        RECT 309.840 59.010 311.050 60.100 ;
        RECT 309.840 58.470 310.360 59.010 ;
        RECT 310.530 58.300 311.050 58.840 ;
        RECT 304.320 57.550 309.665 58.095 ;
        RECT 309.840 57.550 311.050 58.300 ;
        RECT 162.095 57.380 311.135 57.550 ;
        RECT 162.180 56.630 163.390 57.380 ;
        RECT 163.560 56.835 168.905 57.380 ;
        RECT 162.180 56.090 162.700 56.630 ;
        RECT 162.870 55.920 163.390 56.460 ;
        RECT 165.145 56.005 165.485 56.835 ;
        RECT 169.080 56.630 170.290 57.380 ;
        RECT 170.465 56.640 170.720 57.210 ;
        RECT 170.890 56.980 171.220 57.380 ;
        RECT 171.645 56.845 172.175 57.210 ;
        RECT 172.365 57.040 172.640 57.210 ;
        RECT 172.360 56.870 172.640 57.040 ;
        RECT 171.645 56.810 171.820 56.845 ;
        RECT 170.890 56.640 171.820 56.810 ;
        RECT 162.180 54.830 163.390 55.920 ;
        RECT 166.965 55.265 167.315 56.515 ;
        RECT 169.080 56.090 169.600 56.630 ;
        RECT 169.770 55.920 170.290 56.460 ;
        RECT 163.560 54.830 168.905 55.265 ;
        RECT 169.080 54.830 170.290 55.920 ;
        RECT 170.465 55.970 170.635 56.640 ;
        RECT 170.890 56.470 171.060 56.640 ;
        RECT 170.805 56.140 171.060 56.470 ;
        RECT 171.285 56.140 171.480 56.470 ;
        RECT 170.465 55.000 170.800 55.970 ;
        RECT 170.970 54.830 171.140 55.970 ;
        RECT 171.310 55.170 171.480 56.140 ;
        RECT 171.650 55.510 171.820 56.640 ;
        RECT 171.990 55.850 172.160 56.650 ;
        RECT 172.365 56.050 172.640 56.870 ;
        RECT 172.810 55.850 173.000 57.210 ;
        RECT 173.180 56.845 173.690 57.380 ;
        RECT 173.910 56.570 174.155 57.175 ;
        RECT 173.200 56.400 174.430 56.570 ;
        RECT 174.605 56.540 174.865 57.380 ;
        RECT 175.040 56.635 175.295 57.210 ;
        RECT 175.465 57.000 175.795 57.380 ;
        RECT 176.010 56.830 176.180 57.210 ;
        RECT 175.465 56.660 176.180 56.830 ;
        RECT 171.990 55.680 173.000 55.850 ;
        RECT 173.170 55.835 173.920 56.025 ;
        RECT 171.650 55.340 172.775 55.510 ;
        RECT 173.170 55.170 173.340 55.835 ;
        RECT 174.090 55.590 174.430 56.400 ;
        RECT 171.310 55.000 173.340 55.170 ;
        RECT 173.510 54.830 173.680 55.590 ;
        RECT 173.915 55.180 174.430 55.590 ;
        RECT 174.605 54.830 174.865 55.980 ;
        RECT 175.040 55.905 175.210 56.635 ;
        RECT 175.465 56.470 175.635 56.660 ;
        RECT 176.440 56.580 176.730 57.380 ;
        RECT 176.900 56.920 177.450 57.210 ;
        RECT 177.620 56.920 177.870 57.380 ;
        RECT 175.380 56.140 175.635 56.470 ;
        RECT 175.465 55.930 175.635 56.140 ;
        RECT 175.915 56.110 176.270 56.480 ;
        RECT 175.040 55.000 175.295 55.905 ;
        RECT 175.465 55.760 176.180 55.930 ;
        RECT 175.465 54.830 175.795 55.590 ;
        RECT 176.010 55.000 176.180 55.760 ;
        RECT 176.440 54.830 176.730 55.970 ;
        RECT 176.900 55.550 177.150 56.920 ;
        RECT 178.500 56.750 178.830 57.110 ;
        RECT 177.440 56.560 178.830 56.750 ;
        RECT 179.200 56.880 179.500 57.210 ;
        RECT 179.670 56.900 179.945 57.380 ;
        RECT 177.440 56.470 177.610 56.560 ;
        RECT 177.320 56.140 177.610 56.470 ;
        RECT 177.780 56.140 178.110 56.390 ;
        RECT 178.340 56.140 179.030 56.390 ;
        RECT 177.440 55.890 177.610 56.140 ;
        RECT 177.440 55.720 178.380 55.890 ;
        RECT 176.900 55.000 177.350 55.550 ;
        RECT 177.540 54.830 177.870 55.550 ;
        RECT 178.080 55.170 178.380 55.720 ;
        RECT 178.715 55.700 179.030 56.140 ;
        RECT 179.200 55.970 179.370 56.880 ;
        RECT 180.125 56.730 180.420 57.120 ;
        RECT 180.590 56.900 180.845 57.380 ;
        RECT 181.020 56.730 181.280 57.120 ;
        RECT 181.450 56.900 181.730 57.380 ;
        RECT 179.540 56.140 179.890 56.710 ;
        RECT 180.125 56.560 181.775 56.730 ;
        RECT 180.060 56.220 181.200 56.390 ;
        RECT 180.060 55.970 180.230 56.220 ;
        RECT 181.370 56.050 181.775 56.560 ;
        RECT 181.960 56.610 183.630 57.380 ;
        RECT 184.305 56.920 185.055 57.210 ;
        RECT 185.565 56.920 185.895 57.380 ;
        RECT 181.960 56.090 182.710 56.610 ;
        RECT 179.200 55.800 180.230 55.970 ;
        RECT 181.020 55.880 181.775 56.050 ;
        RECT 182.880 55.920 183.630 56.440 ;
        RECT 178.550 54.830 178.830 55.500 ;
        RECT 179.200 55.000 179.510 55.800 ;
        RECT 181.020 55.630 181.280 55.880 ;
        RECT 179.680 54.830 179.990 55.630 ;
        RECT 180.160 55.460 181.280 55.630 ;
        RECT 180.160 55.000 180.420 55.460 ;
        RECT 180.590 54.830 180.845 55.290 ;
        RECT 181.020 55.000 181.280 55.460 ;
        RECT 181.450 54.830 181.735 55.700 ;
        RECT 181.960 54.830 183.630 55.920 ;
        RECT 184.305 55.630 184.675 56.920 ;
        RECT 186.115 56.730 186.385 56.940 ;
        RECT 185.050 56.560 186.385 56.730 ;
        RECT 186.560 56.630 187.770 57.380 ;
        RECT 187.940 56.655 188.230 57.380 ;
        RECT 188.405 57.125 188.740 57.170 ;
        RECT 188.400 56.660 188.740 57.125 ;
        RECT 188.910 57.000 189.240 57.380 ;
        RECT 185.050 56.390 185.220 56.560 ;
        RECT 184.845 56.140 185.220 56.390 ;
        RECT 185.390 56.150 185.865 56.390 ;
        RECT 186.035 56.150 186.385 56.390 ;
        RECT 185.050 55.970 185.220 56.140 ;
        RECT 186.560 56.090 187.080 56.630 ;
        RECT 185.050 55.800 186.385 55.970 ;
        RECT 187.250 55.920 187.770 56.460 ;
        RECT 186.105 55.640 186.385 55.800 ;
        RECT 184.305 55.460 185.475 55.630 ;
        RECT 184.760 54.830 184.975 55.290 ;
        RECT 185.145 55.000 185.475 55.460 ;
        RECT 185.645 54.830 185.895 55.630 ;
        RECT 186.560 54.830 187.770 55.920 ;
        RECT 187.940 54.830 188.230 55.995 ;
        RECT 188.400 55.970 188.570 56.660 ;
        RECT 188.740 56.140 189.000 56.470 ;
        RECT 188.400 55.000 188.660 55.970 ;
        RECT 188.830 55.590 189.000 56.140 ;
        RECT 189.170 55.770 189.510 56.800 ;
        RECT 189.700 56.020 189.970 57.045 ;
        RECT 189.700 55.850 190.010 56.020 ;
        RECT 189.700 55.770 189.970 55.850 ;
        RECT 190.195 55.770 190.475 57.045 ;
        RECT 190.675 56.880 190.905 57.210 ;
        RECT 191.150 57.000 191.480 57.380 ;
        RECT 190.675 55.590 190.845 56.880 ;
        RECT 191.650 56.810 191.825 57.210 ;
        RECT 191.195 56.640 191.825 56.810 ;
        RECT 192.080 56.705 192.340 57.210 ;
        RECT 192.520 57.000 192.850 57.380 ;
        RECT 193.030 56.830 193.200 57.210 ;
        RECT 191.195 56.470 191.365 56.640 ;
        RECT 191.015 56.140 191.365 56.470 ;
        RECT 188.830 55.420 190.845 55.590 ;
        RECT 191.195 55.620 191.365 56.140 ;
        RECT 191.545 55.790 191.910 56.470 ;
        RECT 192.080 55.905 192.260 56.705 ;
        RECT 192.535 56.660 193.200 56.830 ;
        RECT 194.385 56.830 194.640 57.120 ;
        RECT 194.810 57.000 195.140 57.380 ;
        RECT 194.385 56.660 195.135 56.830 ;
        RECT 192.535 56.405 192.705 56.660 ;
        RECT 192.430 56.075 192.705 56.405 ;
        RECT 192.930 56.110 193.270 56.480 ;
        RECT 192.535 55.930 192.705 56.075 ;
        RECT 191.195 55.450 191.825 55.620 ;
        RECT 188.855 54.830 189.185 55.240 ;
        RECT 189.385 55.000 189.555 55.420 ;
        RECT 189.770 54.830 190.440 55.240 ;
        RECT 190.675 55.000 190.845 55.420 ;
        RECT 191.150 54.830 191.480 55.270 ;
        RECT 191.650 55.000 191.825 55.450 ;
        RECT 192.080 55.000 192.350 55.905 ;
        RECT 192.535 55.760 193.210 55.930 ;
        RECT 194.385 55.840 194.735 56.490 ;
        RECT 192.520 54.830 192.850 55.590 ;
        RECT 193.030 55.000 193.210 55.760 ;
        RECT 194.905 55.670 195.135 56.660 ;
        RECT 194.385 55.500 195.135 55.670 ;
        RECT 194.385 55.000 194.640 55.500 ;
        RECT 194.810 54.830 195.140 55.330 ;
        RECT 195.310 55.000 195.480 57.120 ;
        RECT 195.840 57.020 196.170 57.380 ;
        RECT 196.340 56.990 196.835 57.160 ;
        RECT 197.040 56.990 197.895 57.160 ;
        RECT 195.710 55.800 196.170 56.850 ;
        RECT 195.650 55.015 195.975 55.800 ;
        RECT 196.340 55.630 196.510 56.990 ;
        RECT 196.680 56.080 197.030 56.700 ;
        RECT 197.200 56.480 197.555 56.700 ;
        RECT 197.200 55.890 197.370 56.480 ;
        RECT 197.725 56.280 197.895 56.990 ;
        RECT 198.770 56.920 199.100 57.380 ;
        RECT 199.310 57.020 199.660 57.190 ;
        RECT 198.100 56.450 198.890 56.700 ;
        RECT 199.310 56.630 199.570 57.020 ;
        RECT 199.880 56.930 200.830 57.210 ;
        RECT 201.000 56.940 201.190 57.380 ;
        RECT 201.360 57.000 202.430 57.170 ;
        RECT 199.060 56.280 199.230 56.460 ;
        RECT 196.340 55.460 196.735 55.630 ;
        RECT 196.905 55.500 197.370 55.890 ;
        RECT 197.540 56.110 199.230 56.280 ;
        RECT 196.565 55.330 196.735 55.460 ;
        RECT 197.540 55.330 197.710 56.110 ;
        RECT 199.400 55.940 199.570 56.630 ;
        RECT 198.070 55.770 199.570 55.940 ;
        RECT 199.760 55.970 199.970 56.760 ;
        RECT 200.140 56.140 200.490 56.760 ;
        RECT 200.660 56.150 200.830 56.930 ;
        RECT 201.360 56.770 201.530 57.000 ;
        RECT 201.000 56.600 201.530 56.770 ;
        RECT 201.000 56.320 201.220 56.600 ;
        RECT 201.700 56.430 201.940 56.830 ;
        RECT 200.660 55.980 201.065 56.150 ;
        RECT 201.400 56.060 201.940 56.430 ;
        RECT 202.110 56.645 202.430 57.000 ;
        RECT 202.675 56.920 202.980 57.380 ;
        RECT 203.150 56.670 203.405 57.200 ;
        RECT 202.110 56.470 202.435 56.645 ;
        RECT 202.110 56.170 203.025 56.470 ;
        RECT 202.285 56.140 203.025 56.170 ;
        RECT 199.760 55.810 200.435 55.970 ;
        RECT 200.895 55.890 201.065 55.980 ;
        RECT 199.760 55.800 200.725 55.810 ;
        RECT 199.400 55.630 199.570 55.770 ;
        RECT 196.145 54.830 196.395 55.290 ;
        RECT 196.565 55.000 196.815 55.330 ;
        RECT 197.030 55.000 197.710 55.330 ;
        RECT 197.880 55.430 198.955 55.600 ;
        RECT 199.400 55.460 199.960 55.630 ;
        RECT 200.265 55.510 200.725 55.800 ;
        RECT 200.895 55.720 202.115 55.890 ;
        RECT 197.880 55.090 198.050 55.430 ;
        RECT 198.285 54.830 198.615 55.260 ;
        RECT 198.785 55.090 198.955 55.430 ;
        RECT 199.250 54.830 199.620 55.290 ;
        RECT 199.790 55.000 199.960 55.460 ;
        RECT 200.895 55.340 201.065 55.720 ;
        RECT 202.285 55.550 202.455 56.140 ;
        RECT 203.195 56.020 203.405 56.670 ;
        RECT 200.195 55.000 201.065 55.340 ;
        RECT 201.655 55.380 202.455 55.550 ;
        RECT 201.235 54.830 201.485 55.290 ;
        RECT 201.655 55.090 201.825 55.380 ;
        RECT 202.005 54.830 202.335 55.210 ;
        RECT 202.675 54.830 202.980 55.970 ;
        RECT 203.150 55.140 203.405 56.020 ;
        RECT 203.615 56.640 204.230 57.210 ;
        RECT 204.400 56.870 204.615 57.380 ;
        RECT 204.845 56.870 205.125 57.200 ;
        RECT 205.305 56.870 205.545 57.380 ;
        RECT 203.615 55.620 203.930 56.640 ;
        RECT 204.100 55.970 204.270 56.470 ;
        RECT 204.520 56.140 204.785 56.700 ;
        RECT 204.955 55.970 205.125 56.870 ;
        RECT 205.295 56.140 205.650 56.700 ;
        RECT 205.880 56.610 208.470 57.380 ;
        RECT 209.135 56.640 209.750 57.210 ;
        RECT 209.920 56.870 210.135 57.380 ;
        RECT 210.365 56.870 210.645 57.200 ;
        RECT 210.825 56.870 211.065 57.380 ;
        RECT 211.565 56.870 211.805 57.380 ;
        RECT 211.985 56.870 212.265 57.200 ;
        RECT 212.495 56.870 212.710 57.380 ;
        RECT 205.880 56.090 207.090 56.610 ;
        RECT 204.100 55.800 205.525 55.970 ;
        RECT 207.260 55.920 208.470 56.440 ;
        RECT 203.615 55.000 204.150 55.620 ;
        RECT 204.320 54.830 204.650 55.630 ;
        RECT 205.135 55.625 205.525 55.800 ;
        RECT 205.880 54.830 208.470 55.920 ;
        RECT 209.135 55.620 209.450 56.640 ;
        RECT 209.620 55.970 209.790 56.470 ;
        RECT 210.040 56.140 210.305 56.700 ;
        RECT 210.475 55.970 210.645 56.870 ;
        RECT 210.815 56.140 211.170 56.700 ;
        RECT 211.460 56.140 211.815 56.700 ;
        RECT 211.985 55.970 212.155 56.870 ;
        RECT 212.325 56.140 212.590 56.700 ;
        RECT 212.880 56.640 213.495 57.210 ;
        RECT 213.700 56.655 213.990 57.380 ;
        RECT 212.840 55.970 213.010 56.470 ;
        RECT 209.620 55.800 211.045 55.970 ;
        RECT 209.135 55.000 209.670 55.620 ;
        RECT 209.840 54.830 210.170 55.630 ;
        RECT 210.655 55.625 211.045 55.800 ;
        RECT 211.585 55.800 213.010 55.970 ;
        RECT 211.585 55.625 211.975 55.800 ;
        RECT 212.460 54.830 212.790 55.630 ;
        RECT 213.180 55.620 213.495 56.640 ;
        RECT 214.160 56.640 214.600 57.200 ;
        RECT 214.770 56.640 215.220 57.380 ;
        RECT 215.390 56.810 215.560 57.210 ;
        RECT 215.730 56.980 216.150 57.380 ;
        RECT 216.320 56.810 216.550 57.210 ;
        RECT 215.390 56.640 216.550 56.810 ;
        RECT 216.720 56.640 217.210 57.210 ;
        RECT 212.960 55.000 213.495 55.620 ;
        RECT 213.700 54.830 213.990 55.995 ;
        RECT 214.160 55.630 214.470 56.640 ;
        RECT 214.640 56.020 214.810 56.470 ;
        RECT 214.980 56.190 215.370 56.470 ;
        RECT 215.555 56.140 215.800 56.470 ;
        RECT 214.640 55.850 215.430 56.020 ;
        RECT 214.160 55.000 214.600 55.630 ;
        RECT 214.775 54.830 215.090 55.680 ;
        RECT 215.260 55.170 215.430 55.850 ;
        RECT 215.600 55.340 215.800 56.140 ;
        RECT 216.000 55.340 216.250 56.470 ;
        RECT 216.465 56.140 216.870 56.470 ;
        RECT 217.040 55.970 217.210 56.640 ;
        RECT 216.440 55.800 217.210 55.970 ;
        RECT 218.305 56.670 218.560 57.200 ;
        RECT 218.730 56.920 219.035 57.380 ;
        RECT 219.280 57.000 220.350 57.170 ;
        RECT 218.305 56.020 218.515 56.670 ;
        RECT 219.280 56.645 219.600 57.000 ;
        RECT 219.275 56.470 219.600 56.645 ;
        RECT 218.685 56.170 219.600 56.470 ;
        RECT 219.770 56.430 220.010 56.830 ;
        RECT 220.180 56.770 220.350 57.000 ;
        RECT 220.520 56.940 220.710 57.380 ;
        RECT 220.880 56.930 221.830 57.210 ;
        RECT 222.050 57.020 222.400 57.190 ;
        RECT 220.180 56.600 220.710 56.770 ;
        RECT 218.685 56.140 219.425 56.170 ;
        RECT 216.440 55.170 216.690 55.800 ;
        RECT 215.260 55.000 216.690 55.170 ;
        RECT 216.870 54.830 217.200 55.630 ;
        RECT 218.305 55.140 218.560 56.020 ;
        RECT 218.730 54.830 219.035 55.970 ;
        RECT 219.255 55.550 219.425 56.140 ;
        RECT 219.770 56.060 220.310 56.430 ;
        RECT 220.490 56.320 220.710 56.600 ;
        RECT 220.880 56.150 221.050 56.930 ;
        RECT 220.645 55.980 221.050 56.150 ;
        RECT 221.220 56.140 221.570 56.760 ;
        RECT 220.645 55.890 220.815 55.980 ;
        RECT 221.740 55.970 221.950 56.760 ;
        RECT 219.595 55.720 220.815 55.890 ;
        RECT 221.275 55.810 221.950 55.970 ;
        RECT 219.255 55.380 220.055 55.550 ;
        RECT 219.375 54.830 219.705 55.210 ;
        RECT 219.885 55.090 220.055 55.380 ;
        RECT 220.645 55.340 220.815 55.720 ;
        RECT 220.985 55.800 221.950 55.810 ;
        RECT 222.140 56.630 222.400 57.020 ;
        RECT 222.610 56.920 222.940 57.380 ;
        RECT 223.815 56.990 224.670 57.160 ;
        RECT 224.875 56.990 225.370 57.160 ;
        RECT 225.540 57.020 225.870 57.380 ;
        RECT 222.140 55.940 222.310 56.630 ;
        RECT 222.480 56.280 222.650 56.460 ;
        RECT 222.820 56.450 223.610 56.700 ;
        RECT 223.815 56.280 223.985 56.990 ;
        RECT 224.155 56.480 224.510 56.700 ;
        RECT 222.480 56.110 224.170 56.280 ;
        RECT 220.985 55.510 221.445 55.800 ;
        RECT 222.140 55.770 223.640 55.940 ;
        RECT 222.140 55.630 222.310 55.770 ;
        RECT 221.750 55.460 222.310 55.630 ;
        RECT 220.225 54.830 220.475 55.290 ;
        RECT 220.645 55.000 221.515 55.340 ;
        RECT 221.750 55.000 221.920 55.460 ;
        RECT 222.755 55.430 223.830 55.600 ;
        RECT 222.090 54.830 222.460 55.290 ;
        RECT 222.755 55.090 222.925 55.430 ;
        RECT 223.095 54.830 223.425 55.260 ;
        RECT 223.660 55.090 223.830 55.430 ;
        RECT 224.000 55.330 224.170 56.110 ;
        RECT 224.340 55.890 224.510 56.480 ;
        RECT 224.680 56.080 225.030 56.700 ;
        RECT 224.340 55.500 224.805 55.890 ;
        RECT 225.200 55.630 225.370 56.990 ;
        RECT 225.540 55.800 226.000 56.850 ;
        RECT 224.975 55.460 225.370 55.630 ;
        RECT 224.975 55.330 225.145 55.460 ;
        RECT 224.000 55.000 224.680 55.330 ;
        RECT 224.895 55.000 225.145 55.330 ;
        RECT 225.315 54.830 225.565 55.290 ;
        RECT 225.735 55.015 226.060 55.800 ;
        RECT 226.230 55.000 226.400 57.120 ;
        RECT 226.570 57.000 226.900 57.380 ;
        RECT 227.070 56.830 227.325 57.120 ;
        RECT 226.575 56.660 227.325 56.830 ;
        RECT 227.505 56.830 227.760 57.120 ;
        RECT 227.930 57.000 228.260 57.380 ;
        RECT 227.505 56.660 228.255 56.830 ;
        RECT 226.575 55.670 226.805 56.660 ;
        RECT 226.975 55.840 227.325 56.490 ;
        RECT 227.505 55.840 227.855 56.490 ;
        RECT 228.025 55.670 228.255 56.660 ;
        RECT 226.575 55.500 227.325 55.670 ;
        RECT 226.570 54.830 226.900 55.330 ;
        RECT 227.070 55.000 227.325 55.500 ;
        RECT 227.505 55.500 228.255 55.670 ;
        RECT 227.505 55.000 227.760 55.500 ;
        RECT 227.930 54.830 228.260 55.330 ;
        RECT 228.430 55.000 228.600 57.120 ;
        RECT 228.960 57.020 229.290 57.380 ;
        RECT 229.460 56.990 229.955 57.160 ;
        RECT 230.160 56.990 231.015 57.160 ;
        RECT 228.830 55.800 229.290 56.850 ;
        RECT 228.770 55.015 229.095 55.800 ;
        RECT 229.460 55.630 229.630 56.990 ;
        RECT 229.800 56.080 230.150 56.700 ;
        RECT 230.320 56.480 230.675 56.700 ;
        RECT 230.320 55.890 230.490 56.480 ;
        RECT 230.845 56.280 231.015 56.990 ;
        RECT 231.890 56.920 232.220 57.380 ;
        RECT 232.430 57.020 232.780 57.190 ;
        RECT 231.220 56.450 232.010 56.700 ;
        RECT 232.430 56.630 232.690 57.020 ;
        RECT 233.000 56.930 233.950 57.210 ;
        RECT 234.120 56.940 234.310 57.380 ;
        RECT 234.480 57.000 235.550 57.170 ;
        RECT 232.180 56.280 232.350 56.460 ;
        RECT 229.460 55.460 229.855 55.630 ;
        RECT 230.025 55.500 230.490 55.890 ;
        RECT 230.660 56.110 232.350 56.280 ;
        RECT 229.685 55.330 229.855 55.460 ;
        RECT 230.660 55.330 230.830 56.110 ;
        RECT 232.520 55.940 232.690 56.630 ;
        RECT 231.190 55.770 232.690 55.940 ;
        RECT 232.880 55.970 233.090 56.760 ;
        RECT 233.260 56.140 233.610 56.760 ;
        RECT 233.780 56.150 233.950 56.930 ;
        RECT 234.480 56.770 234.650 57.000 ;
        RECT 234.120 56.600 234.650 56.770 ;
        RECT 234.120 56.320 234.340 56.600 ;
        RECT 234.820 56.430 235.060 56.830 ;
        RECT 233.780 55.980 234.185 56.150 ;
        RECT 234.520 56.060 235.060 56.430 ;
        RECT 235.230 56.645 235.550 57.000 ;
        RECT 235.795 56.920 236.100 57.380 ;
        RECT 236.270 56.670 236.525 57.200 ;
        RECT 236.865 56.870 237.105 57.380 ;
        RECT 237.285 56.870 237.565 57.200 ;
        RECT 237.795 56.870 238.010 57.380 ;
        RECT 235.230 56.470 235.555 56.645 ;
        RECT 235.230 56.170 236.145 56.470 ;
        RECT 235.405 56.140 236.145 56.170 ;
        RECT 232.880 55.810 233.555 55.970 ;
        RECT 234.015 55.890 234.185 55.980 ;
        RECT 232.880 55.800 233.845 55.810 ;
        RECT 232.520 55.630 232.690 55.770 ;
        RECT 229.265 54.830 229.515 55.290 ;
        RECT 229.685 55.000 229.935 55.330 ;
        RECT 230.150 55.000 230.830 55.330 ;
        RECT 231.000 55.430 232.075 55.600 ;
        RECT 232.520 55.460 233.080 55.630 ;
        RECT 233.385 55.510 233.845 55.800 ;
        RECT 234.015 55.720 235.235 55.890 ;
        RECT 231.000 55.090 231.170 55.430 ;
        RECT 231.405 54.830 231.735 55.260 ;
        RECT 231.905 55.090 232.075 55.430 ;
        RECT 232.370 54.830 232.740 55.290 ;
        RECT 232.910 55.000 233.080 55.460 ;
        RECT 234.015 55.340 234.185 55.720 ;
        RECT 235.405 55.550 235.575 56.140 ;
        RECT 236.315 56.020 236.525 56.670 ;
        RECT 236.760 56.140 237.115 56.700 ;
        RECT 233.315 55.000 234.185 55.340 ;
        RECT 234.775 55.380 235.575 55.550 ;
        RECT 234.355 54.830 234.605 55.290 ;
        RECT 234.775 55.090 234.945 55.380 ;
        RECT 235.125 54.830 235.455 55.210 ;
        RECT 235.795 54.830 236.100 55.970 ;
        RECT 236.270 55.140 236.525 56.020 ;
        RECT 237.285 55.970 237.455 56.870 ;
        RECT 237.625 56.140 237.890 56.700 ;
        RECT 238.180 56.640 238.795 57.210 ;
        RECT 239.460 56.655 239.750 57.380 ;
        RECT 238.140 55.970 238.310 56.470 ;
        RECT 236.885 55.800 238.310 55.970 ;
        RECT 236.885 55.625 237.275 55.800 ;
        RECT 237.760 54.830 238.090 55.630 ;
        RECT 238.480 55.620 238.795 56.640 ;
        RECT 239.920 56.640 240.305 57.210 ;
        RECT 240.475 56.920 240.800 57.380 ;
        RECT 241.320 56.750 241.600 57.210 ;
        RECT 238.260 55.000 238.795 55.620 ;
        RECT 239.460 54.830 239.750 55.995 ;
        RECT 239.920 55.970 240.200 56.640 ;
        RECT 240.475 56.580 241.600 56.750 ;
        RECT 240.475 56.470 240.925 56.580 ;
        RECT 240.370 56.140 240.925 56.470 ;
        RECT 241.790 56.410 242.190 57.210 ;
        RECT 242.590 56.920 242.860 57.380 ;
        RECT 243.030 56.750 243.315 57.210 ;
        RECT 239.920 55.000 240.305 55.970 ;
        RECT 240.475 55.680 240.925 56.140 ;
        RECT 241.095 55.850 242.190 56.410 ;
        RECT 240.475 55.460 241.600 55.680 ;
        RECT 240.475 54.830 240.800 55.290 ;
        RECT 241.320 55.000 241.600 55.460 ;
        RECT 241.790 55.000 242.190 55.850 ;
        RECT 242.360 56.580 243.315 56.750 ;
        RECT 243.635 56.640 244.250 57.210 ;
        RECT 244.420 56.870 244.635 57.380 ;
        RECT 244.865 56.870 245.145 57.200 ;
        RECT 245.325 56.870 245.565 57.380 ;
        RECT 242.360 55.680 242.570 56.580 ;
        RECT 242.740 55.850 243.430 56.410 ;
        RECT 242.360 55.460 243.315 55.680 ;
        RECT 242.590 54.830 242.860 55.290 ;
        RECT 243.030 55.000 243.315 55.460 ;
        RECT 243.635 55.620 243.950 56.640 ;
        RECT 244.120 55.970 244.290 56.470 ;
        RECT 244.540 56.140 244.805 56.700 ;
        RECT 244.975 55.970 245.145 56.870 ;
        RECT 245.315 56.140 245.670 56.700 ;
        RECT 245.900 56.630 247.110 57.380 ;
        RECT 247.395 56.750 247.680 57.210 ;
        RECT 247.850 56.920 248.120 57.380 ;
        RECT 245.900 56.090 246.420 56.630 ;
        RECT 247.395 56.580 248.350 56.750 ;
        RECT 244.120 55.800 245.545 55.970 ;
        RECT 246.590 55.920 247.110 56.460 ;
        RECT 243.635 55.000 244.170 55.620 ;
        RECT 244.340 54.830 244.670 55.630 ;
        RECT 245.155 55.625 245.545 55.800 ;
        RECT 245.900 54.830 247.110 55.920 ;
        RECT 247.280 55.850 247.970 56.410 ;
        RECT 248.140 55.680 248.350 56.580 ;
        RECT 247.395 55.460 248.350 55.680 ;
        RECT 248.520 56.410 248.920 57.210 ;
        RECT 249.110 56.750 249.390 57.210 ;
        RECT 249.910 56.920 250.235 57.380 ;
        RECT 249.110 56.580 250.235 56.750 ;
        RECT 250.405 56.640 250.790 57.210 ;
        RECT 249.785 56.470 250.235 56.580 ;
        RECT 248.520 55.850 249.615 56.410 ;
        RECT 249.785 56.140 250.340 56.470 ;
        RECT 247.395 55.000 247.680 55.460 ;
        RECT 247.850 54.830 248.120 55.290 ;
        RECT 248.520 55.000 248.920 55.850 ;
        RECT 249.785 55.680 250.235 56.140 ;
        RECT 250.510 55.970 250.790 56.640 ;
        RECT 249.110 55.460 250.235 55.680 ;
        RECT 249.110 55.000 249.390 55.460 ;
        RECT 249.910 54.830 250.235 55.290 ;
        RECT 250.405 55.000 250.790 55.970 ;
        RECT 250.960 56.880 251.220 57.210 ;
        RECT 251.390 57.020 251.720 57.380 ;
        RECT 251.975 57.000 253.275 57.210 ;
        RECT 250.960 55.680 251.130 56.880 ;
        RECT 251.975 56.850 252.145 57.000 ;
        RECT 251.390 56.725 252.145 56.850 ;
        RECT 251.300 56.680 252.145 56.725 ;
        RECT 251.300 56.560 251.570 56.680 ;
        RECT 251.300 55.985 251.470 56.560 ;
        RECT 251.700 56.120 252.110 56.425 ;
        RECT 252.400 56.390 252.610 56.790 ;
        RECT 252.280 56.180 252.610 56.390 ;
        RECT 252.855 56.390 253.075 56.790 ;
        RECT 253.550 56.615 254.005 57.380 ;
        RECT 254.185 56.830 254.440 57.120 ;
        RECT 254.610 57.000 254.940 57.380 ;
        RECT 254.185 56.660 254.935 56.830 ;
        RECT 252.855 56.180 253.330 56.390 ;
        RECT 253.520 56.190 254.010 56.390 ;
        RECT 251.300 55.950 251.500 55.985 ;
        RECT 252.830 55.950 254.005 56.010 ;
        RECT 251.300 55.840 254.005 55.950 ;
        RECT 254.185 55.840 254.535 56.490 ;
        RECT 251.360 55.780 253.160 55.840 ;
        RECT 252.830 55.750 253.160 55.780 ;
        RECT 250.960 55.000 251.220 55.680 ;
        RECT 251.390 54.830 251.640 55.610 ;
        RECT 251.890 55.580 252.725 55.590 ;
        RECT 253.315 55.580 253.500 55.670 ;
        RECT 251.890 55.380 253.500 55.580 ;
        RECT 251.890 55.000 252.140 55.380 ;
        RECT 253.270 55.340 253.500 55.380 ;
        RECT 253.750 55.220 254.005 55.840 ;
        RECT 254.705 55.670 254.935 56.660 ;
        RECT 252.310 54.830 252.665 55.210 ;
        RECT 253.670 55.000 254.005 55.220 ;
        RECT 254.185 55.500 254.935 55.670 ;
        RECT 254.185 55.000 254.440 55.500 ;
        RECT 254.610 54.830 254.940 55.330 ;
        RECT 255.110 55.000 255.280 57.120 ;
        RECT 255.640 57.020 255.970 57.380 ;
        RECT 256.140 56.990 256.635 57.160 ;
        RECT 256.840 56.990 257.695 57.160 ;
        RECT 255.510 55.800 255.970 56.850 ;
        RECT 255.450 55.015 255.775 55.800 ;
        RECT 256.140 55.630 256.310 56.990 ;
        RECT 256.480 56.080 256.830 56.700 ;
        RECT 257.000 56.480 257.355 56.700 ;
        RECT 257.000 55.890 257.170 56.480 ;
        RECT 257.525 56.280 257.695 56.990 ;
        RECT 258.570 56.920 258.900 57.380 ;
        RECT 259.110 57.020 259.460 57.190 ;
        RECT 257.900 56.450 258.690 56.700 ;
        RECT 259.110 56.630 259.370 57.020 ;
        RECT 259.680 56.930 260.630 57.210 ;
        RECT 260.800 56.940 260.990 57.380 ;
        RECT 261.160 57.000 262.230 57.170 ;
        RECT 258.860 56.280 259.030 56.460 ;
        RECT 256.140 55.460 256.535 55.630 ;
        RECT 256.705 55.500 257.170 55.890 ;
        RECT 257.340 56.110 259.030 56.280 ;
        RECT 256.365 55.330 256.535 55.460 ;
        RECT 257.340 55.330 257.510 56.110 ;
        RECT 259.200 55.940 259.370 56.630 ;
        RECT 257.870 55.770 259.370 55.940 ;
        RECT 259.560 55.970 259.770 56.760 ;
        RECT 259.940 56.140 260.290 56.760 ;
        RECT 260.460 56.150 260.630 56.930 ;
        RECT 261.160 56.770 261.330 57.000 ;
        RECT 260.800 56.600 261.330 56.770 ;
        RECT 260.800 56.320 261.020 56.600 ;
        RECT 261.500 56.430 261.740 56.830 ;
        RECT 260.460 55.980 260.865 56.150 ;
        RECT 261.200 56.060 261.740 56.430 ;
        RECT 261.910 56.645 262.230 57.000 ;
        RECT 262.475 56.920 262.780 57.380 ;
        RECT 262.950 56.670 263.205 57.200 ;
        RECT 261.910 56.470 262.235 56.645 ;
        RECT 261.910 56.170 262.825 56.470 ;
        RECT 262.085 56.140 262.825 56.170 ;
        RECT 259.560 55.810 260.235 55.970 ;
        RECT 260.695 55.890 260.865 55.980 ;
        RECT 259.560 55.800 260.525 55.810 ;
        RECT 259.200 55.630 259.370 55.770 ;
        RECT 255.945 54.830 256.195 55.290 ;
        RECT 256.365 55.000 256.615 55.330 ;
        RECT 256.830 55.000 257.510 55.330 ;
        RECT 257.680 55.430 258.755 55.600 ;
        RECT 259.200 55.460 259.760 55.630 ;
        RECT 260.065 55.510 260.525 55.800 ;
        RECT 260.695 55.720 261.915 55.890 ;
        RECT 257.680 55.090 257.850 55.430 ;
        RECT 258.085 54.830 258.415 55.260 ;
        RECT 258.585 55.090 258.755 55.430 ;
        RECT 259.050 54.830 259.420 55.290 ;
        RECT 259.590 55.000 259.760 55.460 ;
        RECT 260.695 55.340 260.865 55.720 ;
        RECT 262.085 55.550 262.255 56.140 ;
        RECT 262.995 56.020 263.205 56.670 ;
        RECT 263.420 56.560 263.650 57.380 ;
        RECT 263.820 56.580 264.150 57.210 ;
        RECT 263.400 56.140 263.730 56.390 ;
        RECT 259.995 55.000 260.865 55.340 ;
        RECT 261.455 55.380 262.255 55.550 ;
        RECT 261.035 54.830 261.285 55.290 ;
        RECT 261.455 55.090 261.625 55.380 ;
        RECT 261.805 54.830 262.135 55.210 ;
        RECT 262.475 54.830 262.780 55.970 ;
        RECT 262.950 55.140 263.205 56.020 ;
        RECT 263.900 55.980 264.150 56.580 ;
        RECT 264.320 56.560 264.530 57.380 ;
        RECT 265.220 56.655 265.510 57.380 ;
        RECT 265.680 56.835 271.025 57.380 ;
        RECT 267.265 56.005 267.605 56.835 ;
        RECT 271.200 56.610 274.710 57.380 ;
        RECT 275.345 56.830 275.600 57.120 ;
        RECT 275.770 57.000 276.100 57.380 ;
        RECT 275.345 56.660 276.095 56.830 ;
        RECT 263.420 54.830 263.650 55.970 ;
        RECT 263.820 55.000 264.150 55.980 ;
        RECT 264.320 54.830 264.530 55.970 ;
        RECT 265.220 54.830 265.510 55.995 ;
        RECT 269.085 55.265 269.435 56.515 ;
        RECT 271.200 56.090 272.850 56.610 ;
        RECT 273.020 55.920 274.710 56.440 ;
        RECT 265.680 54.830 271.025 55.265 ;
        RECT 271.200 54.830 274.710 55.920 ;
        RECT 275.345 55.840 275.695 56.490 ;
        RECT 275.865 55.670 276.095 56.660 ;
        RECT 275.345 55.500 276.095 55.670 ;
        RECT 275.345 55.000 275.600 55.500 ;
        RECT 275.770 54.830 276.100 55.330 ;
        RECT 276.270 55.000 276.440 57.120 ;
        RECT 276.800 57.020 277.130 57.380 ;
        RECT 277.300 56.990 277.795 57.160 ;
        RECT 278.000 56.990 278.855 57.160 ;
        RECT 276.670 55.800 277.130 56.850 ;
        RECT 276.610 55.015 276.935 55.800 ;
        RECT 277.300 55.630 277.470 56.990 ;
        RECT 277.640 56.080 277.990 56.700 ;
        RECT 278.160 56.480 278.515 56.700 ;
        RECT 278.160 55.890 278.330 56.480 ;
        RECT 278.685 56.280 278.855 56.990 ;
        RECT 279.730 56.920 280.060 57.380 ;
        RECT 280.270 57.020 280.620 57.190 ;
        RECT 279.060 56.450 279.850 56.700 ;
        RECT 280.270 56.630 280.530 57.020 ;
        RECT 280.840 56.930 281.790 57.210 ;
        RECT 281.960 56.940 282.150 57.380 ;
        RECT 282.320 57.000 283.390 57.170 ;
        RECT 280.020 56.280 280.190 56.460 ;
        RECT 277.300 55.460 277.695 55.630 ;
        RECT 277.865 55.500 278.330 55.890 ;
        RECT 278.500 56.110 280.190 56.280 ;
        RECT 277.525 55.330 277.695 55.460 ;
        RECT 278.500 55.330 278.670 56.110 ;
        RECT 280.360 55.940 280.530 56.630 ;
        RECT 279.030 55.770 280.530 55.940 ;
        RECT 280.720 55.970 280.930 56.760 ;
        RECT 281.100 56.140 281.450 56.760 ;
        RECT 281.620 56.150 281.790 56.930 ;
        RECT 282.320 56.770 282.490 57.000 ;
        RECT 281.960 56.600 282.490 56.770 ;
        RECT 281.960 56.320 282.180 56.600 ;
        RECT 282.660 56.430 282.900 56.830 ;
        RECT 281.620 55.980 282.025 56.150 ;
        RECT 282.360 56.060 282.900 56.430 ;
        RECT 283.070 56.645 283.390 57.000 ;
        RECT 283.635 56.920 283.940 57.380 ;
        RECT 284.110 56.670 284.365 57.200 ;
        RECT 284.785 56.900 285.085 57.380 ;
        RECT 285.255 56.730 285.515 57.185 ;
        RECT 285.685 56.900 285.945 57.380 ;
        RECT 286.115 56.730 286.375 57.185 ;
        RECT 286.545 56.900 286.805 57.380 ;
        RECT 286.975 56.730 287.235 57.185 ;
        RECT 287.405 56.900 287.665 57.380 ;
        RECT 287.835 56.730 288.095 57.185 ;
        RECT 288.265 56.855 288.525 57.380 ;
        RECT 283.070 56.470 283.395 56.645 ;
        RECT 283.070 56.170 283.985 56.470 ;
        RECT 283.245 56.140 283.985 56.170 ;
        RECT 280.720 55.810 281.395 55.970 ;
        RECT 281.855 55.890 282.025 55.980 ;
        RECT 280.720 55.800 281.685 55.810 ;
        RECT 280.360 55.630 280.530 55.770 ;
        RECT 277.105 54.830 277.355 55.290 ;
        RECT 277.525 55.000 277.775 55.330 ;
        RECT 277.990 55.000 278.670 55.330 ;
        RECT 278.840 55.430 279.915 55.600 ;
        RECT 280.360 55.460 280.920 55.630 ;
        RECT 281.225 55.510 281.685 55.800 ;
        RECT 281.855 55.720 283.075 55.890 ;
        RECT 278.840 55.090 279.010 55.430 ;
        RECT 279.245 54.830 279.575 55.260 ;
        RECT 279.745 55.090 279.915 55.430 ;
        RECT 280.210 54.830 280.580 55.290 ;
        RECT 280.750 55.000 280.920 55.460 ;
        RECT 281.855 55.340 282.025 55.720 ;
        RECT 283.245 55.550 283.415 56.140 ;
        RECT 284.155 56.020 284.365 56.670 ;
        RECT 281.155 55.000 282.025 55.340 ;
        RECT 282.615 55.380 283.415 55.550 ;
        RECT 282.195 54.830 282.445 55.290 ;
        RECT 282.615 55.090 282.785 55.380 ;
        RECT 282.965 54.830 283.295 55.210 ;
        RECT 283.635 54.830 283.940 55.970 ;
        RECT 284.110 55.140 284.365 56.020 ;
        RECT 284.785 56.560 288.095 56.730 ;
        RECT 284.785 55.970 285.755 56.560 ;
        RECT 288.695 56.390 288.945 57.200 ;
        RECT 289.125 56.920 289.370 57.380 ;
        RECT 285.925 56.140 288.945 56.390 ;
        RECT 289.115 56.140 289.430 56.750 ;
        RECT 289.600 56.630 290.810 57.380 ;
        RECT 290.980 56.655 291.270 57.380 ;
        RECT 291.445 56.640 291.700 57.210 ;
        RECT 291.870 56.980 292.200 57.380 ;
        RECT 292.625 56.845 293.155 57.210 ;
        RECT 293.345 57.040 293.620 57.210 ;
        RECT 293.340 56.870 293.620 57.040 ;
        RECT 292.625 56.810 292.800 56.845 ;
        RECT 291.870 56.640 292.800 56.810 ;
        RECT 284.785 55.730 288.095 55.970 ;
        RECT 284.790 54.830 285.085 55.560 ;
        RECT 285.255 55.005 285.515 55.730 ;
        RECT 285.685 54.830 285.945 55.560 ;
        RECT 286.115 55.005 286.375 55.730 ;
        RECT 286.545 54.830 286.805 55.560 ;
        RECT 286.975 55.005 287.235 55.730 ;
        RECT 287.405 54.830 287.665 55.560 ;
        RECT 287.835 55.005 288.095 55.730 ;
        RECT 288.265 54.830 288.525 55.940 ;
        RECT 288.695 55.005 288.945 56.140 ;
        RECT 289.600 56.090 290.120 56.630 ;
        RECT 289.125 54.830 289.420 55.940 ;
        RECT 290.290 55.920 290.810 56.460 ;
        RECT 289.600 54.830 290.810 55.920 ;
        RECT 290.980 54.830 291.270 55.995 ;
        RECT 291.445 55.970 291.615 56.640 ;
        RECT 291.870 56.470 292.040 56.640 ;
        RECT 291.785 56.140 292.040 56.470 ;
        RECT 292.265 56.140 292.460 56.470 ;
        RECT 291.445 55.000 291.780 55.970 ;
        RECT 291.950 54.830 292.120 55.970 ;
        RECT 292.290 55.170 292.460 56.140 ;
        RECT 292.630 55.510 292.800 56.640 ;
        RECT 292.970 55.850 293.140 56.650 ;
        RECT 293.345 56.050 293.620 56.870 ;
        RECT 293.790 55.850 293.980 57.210 ;
        RECT 294.160 56.845 294.670 57.380 ;
        RECT 294.890 56.570 295.135 57.175 ;
        RECT 295.580 56.610 299.090 57.380 ;
        RECT 299.720 56.870 299.990 57.380 ;
        RECT 300.160 56.700 300.405 57.200 ;
        RECT 299.720 56.640 300.405 56.700 ;
        RECT 300.575 56.640 300.905 57.380 ;
        RECT 299.720 56.610 300.320 56.640 ;
        RECT 294.180 56.400 295.410 56.570 ;
        RECT 292.970 55.680 293.980 55.850 ;
        RECT 294.150 55.835 294.900 56.025 ;
        RECT 292.630 55.340 293.755 55.510 ;
        RECT 294.150 55.170 294.320 55.835 ;
        RECT 295.070 55.590 295.410 56.400 ;
        RECT 295.580 56.090 297.230 56.610 ;
        RECT 299.720 56.570 300.305 56.610 ;
        RECT 297.400 55.920 299.090 56.440 ;
        RECT 292.290 55.000 294.320 55.170 ;
        RECT 294.490 54.830 294.660 55.590 ;
        RECT 294.895 55.180 295.410 55.590 ;
        RECT 295.580 54.830 299.090 55.920 ;
        RECT 299.720 56.020 300.275 56.570 ;
        RECT 301.075 56.470 301.245 57.120 ;
        RECT 300.445 56.140 301.245 56.470 ;
        RECT 299.720 55.970 300.320 56.020 ;
        RECT 299.720 55.850 300.485 55.970 ;
        RECT 299.720 54.830 299.985 55.680 ;
        RECT 300.155 55.005 300.485 55.850 ;
        RECT 300.655 54.830 300.825 55.970 ;
        RECT 300.995 55.550 301.245 56.140 ;
        RECT 301.415 56.785 301.765 57.115 ;
        RECT 301.965 56.900 302.605 57.380 ;
        RECT 302.805 56.990 303.655 57.160 ;
        RECT 301.415 55.890 301.605 56.785 ;
        RECT 301.955 56.460 302.635 56.730 ;
        RECT 302.285 56.400 302.635 56.460 ;
        RECT 301.805 56.230 302.155 56.290 ;
        RECT 302.805 56.230 302.975 56.990 ;
        RECT 304.215 56.920 304.535 57.380 ;
        RECT 304.735 56.740 304.985 57.170 ;
        RECT 305.275 56.940 305.685 57.380 ;
        RECT 305.855 57.000 306.870 57.200 ;
        RECT 303.145 56.570 304.415 56.740 ;
        RECT 303.145 56.450 303.495 56.570 ;
        RECT 301.805 56.060 303.725 56.230 ;
        RECT 301.415 55.720 303.385 55.890 ;
        RECT 301.415 55.700 301.785 55.720 ;
        RECT 300.995 55.040 301.325 55.550 ;
        RECT 301.615 55.090 301.785 55.700 ;
        RECT 303.555 55.550 303.725 56.060 ;
        RECT 303.895 55.990 304.075 56.400 ;
        RECT 304.245 55.810 304.415 56.570 ;
        RECT 301.955 54.830 302.285 55.520 ;
        RECT 302.515 55.380 303.725 55.550 ;
        RECT 303.895 55.500 304.415 55.810 ;
        RECT 304.585 56.400 304.985 56.740 ;
        RECT 305.275 56.400 305.685 56.730 ;
        RECT 304.585 55.630 304.755 56.400 ;
        RECT 305.855 56.270 306.025 57.000 ;
        RECT 307.170 56.830 307.340 57.160 ;
        RECT 307.510 57.000 307.840 57.380 ;
        RECT 308.060 56.900 308.280 57.120 ;
        RECT 308.450 57.000 308.780 57.380 ;
        RECT 306.195 56.450 306.545 56.820 ;
        RECT 305.855 56.230 306.275 56.270 ;
        RECT 304.925 56.060 306.275 56.230 ;
        RECT 304.925 55.900 305.175 56.060 ;
        RECT 305.685 55.630 305.935 55.890 ;
        RECT 304.585 55.380 305.935 55.630 ;
        RECT 302.515 55.090 302.755 55.380 ;
        RECT 303.555 55.300 303.725 55.380 ;
        RECT 302.955 54.830 303.375 55.210 ;
        RECT 303.555 55.050 304.185 55.300 ;
        RECT 304.635 54.830 304.965 55.210 ;
        RECT 305.135 55.090 305.305 55.380 ;
        RECT 306.105 55.215 306.275 56.060 ;
        RECT 306.725 55.890 306.945 56.760 ;
        RECT 307.170 56.640 307.865 56.830 ;
        RECT 306.445 55.510 306.945 55.890 ;
        RECT 307.115 55.840 307.525 56.460 ;
        RECT 307.695 55.670 307.865 56.640 ;
        RECT 307.170 55.500 307.865 55.670 ;
        RECT 305.485 54.830 305.865 55.210 ;
        RECT 306.105 55.045 306.935 55.215 ;
        RECT 307.170 55.000 307.340 55.500 ;
        RECT 308.060 55.420 308.290 56.900 ;
        RECT 308.950 56.830 309.210 57.120 ;
        RECT 308.460 56.660 309.210 56.830 ;
        RECT 308.460 55.670 308.690 56.660 ;
        RECT 309.840 56.630 311.050 57.380 ;
        RECT 308.860 55.840 309.210 56.490 ;
        RECT 309.840 55.920 310.360 56.460 ;
        RECT 310.530 56.090 311.050 56.630 ;
        RECT 308.460 55.500 309.210 55.670 ;
        RECT 307.510 54.830 307.840 55.330 ;
        RECT 308.060 55.000 308.280 55.420 ;
        RECT 308.450 54.830 308.780 55.330 ;
        RECT 308.950 55.000 309.210 55.500 ;
        RECT 309.840 54.830 311.050 55.920 ;
        RECT 162.095 54.660 311.135 54.830 ;
        RECT 162.180 53.570 163.390 54.660 ;
        RECT 163.560 53.570 165.230 54.660 ;
        RECT 165.865 53.990 166.120 54.490 ;
        RECT 166.290 54.160 166.620 54.660 ;
        RECT 165.865 53.820 166.615 53.990 ;
        RECT 162.180 52.860 162.700 53.400 ;
        RECT 162.870 53.030 163.390 53.570 ;
        RECT 163.560 52.880 164.310 53.400 ;
        RECT 164.480 53.050 165.230 53.570 ;
        RECT 165.865 53.000 166.215 53.650 ;
        RECT 162.180 52.110 163.390 52.860 ;
        RECT 163.560 52.110 165.230 52.880 ;
        RECT 166.385 52.830 166.615 53.820 ;
        RECT 165.865 52.660 166.615 52.830 ;
        RECT 165.865 52.370 166.120 52.660 ;
        RECT 166.290 52.110 166.620 52.490 ;
        RECT 166.790 52.370 166.960 54.490 ;
        RECT 167.130 53.690 167.455 54.475 ;
        RECT 167.625 54.200 167.875 54.660 ;
        RECT 168.045 54.160 168.295 54.490 ;
        RECT 168.510 54.160 169.190 54.490 ;
        RECT 168.045 54.030 168.215 54.160 ;
        RECT 167.820 53.860 168.215 54.030 ;
        RECT 167.190 52.640 167.650 53.690 ;
        RECT 167.820 52.500 167.990 53.860 ;
        RECT 168.385 53.600 168.850 53.990 ;
        RECT 168.160 52.790 168.510 53.410 ;
        RECT 168.680 53.010 168.850 53.600 ;
        RECT 169.020 53.380 169.190 54.160 ;
        RECT 169.360 54.060 169.530 54.400 ;
        RECT 169.765 54.230 170.095 54.660 ;
        RECT 170.265 54.060 170.435 54.400 ;
        RECT 170.730 54.200 171.100 54.660 ;
        RECT 169.360 53.890 170.435 54.060 ;
        RECT 171.270 54.030 171.440 54.490 ;
        RECT 171.675 54.150 172.545 54.490 ;
        RECT 172.715 54.200 172.965 54.660 ;
        RECT 170.880 53.860 171.440 54.030 ;
        RECT 170.880 53.720 171.050 53.860 ;
        RECT 169.550 53.550 171.050 53.720 ;
        RECT 171.745 53.690 172.205 53.980 ;
        RECT 169.020 53.210 170.710 53.380 ;
        RECT 168.680 52.790 169.035 53.010 ;
        RECT 169.205 52.500 169.375 53.210 ;
        RECT 169.580 52.790 170.370 53.040 ;
        RECT 170.540 53.030 170.710 53.210 ;
        RECT 170.880 52.860 171.050 53.550 ;
        RECT 167.320 52.110 167.650 52.470 ;
        RECT 167.820 52.330 168.315 52.500 ;
        RECT 168.520 52.330 169.375 52.500 ;
        RECT 170.250 52.110 170.580 52.570 ;
        RECT 170.790 52.470 171.050 52.860 ;
        RECT 171.240 53.680 172.205 53.690 ;
        RECT 172.375 53.770 172.545 54.150 ;
        RECT 173.135 54.110 173.305 54.400 ;
        RECT 173.485 54.280 173.815 54.660 ;
        RECT 173.135 53.940 173.935 54.110 ;
        RECT 171.240 53.520 171.915 53.680 ;
        RECT 172.375 53.600 173.595 53.770 ;
        RECT 171.240 52.730 171.450 53.520 ;
        RECT 172.375 53.510 172.545 53.600 ;
        RECT 171.620 52.730 171.970 53.350 ;
        RECT 172.140 53.340 172.545 53.510 ;
        RECT 172.140 52.560 172.310 53.340 ;
        RECT 172.480 52.890 172.700 53.170 ;
        RECT 172.880 53.060 173.420 53.430 ;
        RECT 173.765 53.350 173.935 53.940 ;
        RECT 174.155 53.520 174.460 54.660 ;
        RECT 174.630 53.470 174.885 54.350 ;
        RECT 175.060 53.495 175.350 54.660 ;
        RECT 175.525 53.520 175.860 54.490 ;
        RECT 176.030 53.520 176.200 54.660 ;
        RECT 176.370 54.320 178.400 54.490 ;
        RECT 173.765 53.320 174.505 53.350 ;
        RECT 172.480 52.720 173.010 52.890 ;
        RECT 170.790 52.300 171.140 52.470 ;
        RECT 171.360 52.280 172.310 52.560 ;
        RECT 172.480 52.110 172.670 52.550 ;
        RECT 172.840 52.490 173.010 52.720 ;
        RECT 173.180 52.660 173.420 53.060 ;
        RECT 173.590 53.020 174.505 53.320 ;
        RECT 173.590 52.845 173.915 53.020 ;
        RECT 173.590 52.490 173.910 52.845 ;
        RECT 174.675 52.820 174.885 53.470 ;
        RECT 175.525 52.850 175.695 53.520 ;
        RECT 176.370 53.350 176.540 54.320 ;
        RECT 175.865 53.020 176.120 53.350 ;
        RECT 176.345 53.020 176.540 53.350 ;
        RECT 176.710 53.980 177.835 54.150 ;
        RECT 175.950 52.850 176.120 53.020 ;
        RECT 176.710 52.850 176.880 53.980 ;
        RECT 172.840 52.320 173.910 52.490 ;
        RECT 174.155 52.110 174.460 52.570 ;
        RECT 174.630 52.290 174.885 52.820 ;
        RECT 175.060 52.110 175.350 52.835 ;
        RECT 175.525 52.280 175.780 52.850 ;
        RECT 175.950 52.680 176.880 52.850 ;
        RECT 177.050 53.640 178.060 53.810 ;
        RECT 177.050 52.840 177.220 53.640 ;
        RECT 177.425 52.960 177.700 53.440 ;
        RECT 177.420 52.790 177.700 52.960 ;
        RECT 176.705 52.645 176.880 52.680 ;
        RECT 175.950 52.110 176.280 52.510 ;
        RECT 176.705 52.280 177.235 52.645 ;
        RECT 177.425 52.280 177.700 52.790 ;
        RECT 177.870 52.280 178.060 53.640 ;
        RECT 178.230 53.655 178.400 54.320 ;
        RECT 178.570 53.900 178.740 54.660 ;
        RECT 178.975 53.900 179.490 54.310 ;
        RECT 178.230 53.465 178.980 53.655 ;
        RECT 179.150 53.090 179.490 53.900 ;
        RECT 179.715 53.790 180.000 54.660 ;
        RECT 180.170 54.030 180.430 54.490 ;
        RECT 180.605 54.200 180.860 54.660 ;
        RECT 181.030 54.030 181.290 54.490 ;
        RECT 180.170 53.860 181.290 54.030 ;
        RECT 181.460 53.860 181.770 54.660 ;
        RECT 180.170 53.610 180.430 53.860 ;
        RECT 181.940 53.690 182.250 54.490 ;
        RECT 182.885 54.280 183.220 54.660 ;
        RECT 178.260 52.920 179.490 53.090 ;
        RECT 179.675 53.440 180.430 53.610 ;
        RECT 181.220 53.520 182.250 53.690 ;
        RECT 179.675 52.930 180.080 53.440 ;
        RECT 181.220 53.270 181.390 53.520 ;
        RECT 180.250 53.100 181.390 53.270 ;
        RECT 178.240 52.110 178.750 52.645 ;
        RECT 178.970 52.315 179.215 52.920 ;
        RECT 179.675 52.760 181.325 52.930 ;
        RECT 181.560 52.780 181.910 53.350 ;
        RECT 179.720 52.110 180.000 52.590 ;
        RECT 180.170 52.370 180.430 52.760 ;
        RECT 180.605 52.110 180.860 52.590 ;
        RECT 181.030 52.370 181.325 52.760 ;
        RECT 182.080 52.610 182.250 53.520 ;
        RECT 182.880 52.790 183.120 54.100 ;
        RECT 183.390 53.690 183.640 54.490 ;
        RECT 183.860 53.940 184.190 54.660 ;
        RECT 184.375 53.690 184.625 54.490 ;
        RECT 185.090 53.860 185.420 54.660 ;
        RECT 185.590 54.230 185.930 54.490 ;
        RECT 183.290 53.520 185.480 53.690 ;
        RECT 183.290 52.610 183.460 53.520 ;
        RECT 185.165 53.350 185.480 53.520 ;
        RECT 181.505 52.110 181.780 52.590 ;
        RECT 181.950 52.280 182.250 52.610 ;
        RECT 182.965 52.280 183.460 52.610 ;
        RECT 183.680 52.385 184.030 53.350 ;
        RECT 184.210 52.380 184.510 53.350 ;
        RECT 184.690 52.380 184.970 53.350 ;
        RECT 185.165 53.100 185.495 53.350 ;
        RECT 185.150 52.110 185.420 52.910 ;
        RECT 185.670 52.830 185.930 54.230 ;
        RECT 186.100 54.150 186.360 54.660 ;
        RECT 186.100 53.100 186.440 53.980 ;
        RECT 186.610 53.270 186.780 54.490 ;
        RECT 187.020 54.155 187.635 54.660 ;
        RECT 187.020 53.620 187.270 53.985 ;
        RECT 187.440 53.980 187.635 54.155 ;
        RECT 187.805 54.150 188.280 54.490 ;
        RECT 188.450 54.115 188.665 54.660 ;
        RECT 187.440 53.790 187.770 53.980 ;
        RECT 187.990 53.620 188.705 53.915 ;
        RECT 188.875 53.790 189.150 54.490 ;
        RECT 190.080 54.020 190.410 54.450 ;
        RECT 187.020 53.450 188.810 53.620 ;
        RECT 186.610 53.020 187.405 53.270 ;
        RECT 186.610 52.930 186.860 53.020 ;
        RECT 185.590 52.320 185.930 52.830 ;
        RECT 186.100 52.110 186.360 52.930 ;
        RECT 186.530 52.510 186.860 52.930 ;
        RECT 187.575 52.595 187.830 53.450 ;
        RECT 187.040 52.330 187.830 52.595 ;
        RECT 188.000 52.750 188.410 53.270 ;
        RECT 188.580 53.020 188.810 53.450 ;
        RECT 188.980 52.760 189.150 53.790 ;
        RECT 188.000 52.330 188.200 52.750 ;
        RECT 188.390 52.110 188.720 52.570 ;
        RECT 188.890 52.280 189.150 52.760 ;
        RECT 189.955 53.850 190.410 54.020 ;
        RECT 190.590 54.020 190.840 54.440 ;
        RECT 191.070 54.190 191.400 54.660 ;
        RECT 191.630 54.020 191.880 54.440 ;
        RECT 190.590 53.850 191.880 54.020 ;
        RECT 189.955 52.850 190.125 53.850 ;
        RECT 190.295 53.020 190.540 53.680 ;
        RECT 190.755 53.020 191.020 53.680 ;
        RECT 191.215 53.020 191.500 53.680 ;
        RECT 191.675 53.350 191.890 53.680 ;
        RECT 192.070 53.520 192.320 54.660 ;
        RECT 192.490 53.600 192.820 54.450 ;
        RECT 193.250 53.930 193.545 54.660 ;
        RECT 193.715 53.760 193.975 54.485 ;
        RECT 194.145 53.930 194.405 54.660 ;
        RECT 194.575 53.760 194.835 54.485 ;
        RECT 195.005 53.930 195.265 54.660 ;
        RECT 195.435 53.760 195.695 54.485 ;
        RECT 195.865 53.930 196.125 54.660 ;
        RECT 196.295 53.760 196.555 54.485 ;
        RECT 192.600 53.470 192.820 53.600 ;
        RECT 191.675 53.020 191.980 53.350 ;
        RECT 192.150 53.020 192.460 53.350 ;
        RECT 192.150 52.850 192.320 53.020 ;
        RECT 189.955 52.680 192.320 52.850 ;
        RECT 192.630 52.835 192.820 53.470 ;
        RECT 190.110 52.110 190.440 52.510 ;
        RECT 190.610 52.340 190.940 52.680 ;
        RECT 191.990 52.110 192.320 52.510 ;
        RECT 192.490 52.325 192.820 52.835 ;
        RECT 193.245 53.520 196.555 53.760 ;
        RECT 196.725 53.550 196.985 54.660 ;
        RECT 193.245 52.930 194.215 53.520 ;
        RECT 197.155 53.350 197.405 54.485 ;
        RECT 197.585 53.550 197.880 54.660 ;
        RECT 198.060 53.520 198.320 54.660 ;
        RECT 198.490 53.690 198.820 54.490 ;
        RECT 198.990 53.860 199.160 54.660 ;
        RECT 199.330 53.690 199.660 54.490 ;
        RECT 199.830 53.860 200.085 54.660 ;
        RECT 198.490 53.520 200.190 53.690 ;
        RECT 194.385 53.100 197.405 53.350 ;
        RECT 193.245 52.760 196.555 52.930 ;
        RECT 193.245 52.110 193.545 52.590 ;
        RECT 193.715 52.305 193.975 52.760 ;
        RECT 194.145 52.110 194.405 52.590 ;
        RECT 194.575 52.305 194.835 52.760 ;
        RECT 195.005 52.110 195.265 52.590 ;
        RECT 195.435 52.305 195.695 52.760 ;
        RECT 195.865 52.110 196.125 52.590 ;
        RECT 196.295 52.305 196.555 52.760 ;
        RECT 196.725 52.110 196.985 52.635 ;
        RECT 197.155 52.290 197.405 53.100 ;
        RECT 197.575 52.740 197.890 53.350 ;
        RECT 198.060 53.100 198.820 53.350 ;
        RECT 198.990 53.100 199.740 53.350 ;
        RECT 199.910 52.930 200.190 53.520 ;
        RECT 200.820 53.495 201.110 54.660 ;
        RECT 201.280 53.570 202.490 54.660 ;
        RECT 198.060 52.740 199.160 52.910 ;
        RECT 197.585 52.110 197.830 52.570 ;
        RECT 198.060 52.280 198.400 52.740 ;
        RECT 198.570 52.110 198.740 52.570 ;
        RECT 198.910 52.490 199.160 52.740 ;
        RECT 199.330 52.680 200.190 52.930 ;
        RECT 201.280 52.860 201.800 53.400 ;
        RECT 201.970 53.030 202.490 53.570 ;
        RECT 202.695 53.870 203.230 54.490 ;
        RECT 199.750 52.490 200.080 52.510 ;
        RECT 198.910 52.280 200.080 52.490 ;
        RECT 200.820 52.110 201.110 52.835 ;
        RECT 201.280 52.110 202.490 52.860 ;
        RECT 202.695 52.850 203.010 53.870 ;
        RECT 203.400 53.860 203.730 54.660 ;
        RECT 205.160 53.990 205.440 54.660 ;
        RECT 204.215 53.690 204.605 53.865 ;
        RECT 205.610 53.770 205.910 54.320 ;
        RECT 206.110 53.940 206.440 54.660 ;
        RECT 206.630 53.940 207.090 54.490 ;
        RECT 203.180 53.520 204.605 53.690 ;
        RECT 203.180 53.020 203.350 53.520 ;
        RECT 202.695 52.280 203.310 52.850 ;
        RECT 203.600 52.790 203.865 53.350 ;
        RECT 204.035 52.620 204.205 53.520 ;
        RECT 204.975 53.350 205.240 53.710 ;
        RECT 205.610 53.600 206.550 53.770 ;
        RECT 206.380 53.350 206.550 53.600 ;
        RECT 204.375 52.790 204.730 53.350 ;
        RECT 204.975 53.100 205.650 53.350 ;
        RECT 205.870 53.100 206.210 53.350 ;
        RECT 206.380 53.020 206.670 53.350 ;
        RECT 206.380 52.930 206.550 53.020 ;
        RECT 205.160 52.740 206.550 52.930 ;
        RECT 203.480 52.110 203.695 52.620 ;
        RECT 203.925 52.290 204.205 52.620 ;
        RECT 204.385 52.110 204.625 52.620 ;
        RECT 205.160 52.380 205.490 52.740 ;
        RECT 206.840 52.570 207.090 53.940 ;
        RECT 207.260 53.570 209.850 54.660 ;
        RECT 210.025 53.990 210.280 54.490 ;
        RECT 210.450 54.160 210.780 54.660 ;
        RECT 210.025 53.820 210.775 53.990 ;
        RECT 206.110 52.110 206.360 52.570 ;
        RECT 206.530 52.280 207.090 52.570 ;
        RECT 207.260 52.880 208.470 53.400 ;
        RECT 208.640 53.050 209.850 53.570 ;
        RECT 210.025 53.000 210.375 53.650 ;
        RECT 207.260 52.110 209.850 52.880 ;
        RECT 210.545 52.830 210.775 53.820 ;
        RECT 210.025 52.660 210.775 52.830 ;
        RECT 210.025 52.370 210.280 52.660 ;
        RECT 210.450 52.110 210.780 52.490 ;
        RECT 210.950 52.370 211.120 54.490 ;
        RECT 211.290 53.690 211.615 54.475 ;
        RECT 211.785 54.200 212.035 54.660 ;
        RECT 212.205 54.160 212.455 54.490 ;
        RECT 212.670 54.160 213.350 54.490 ;
        RECT 212.205 54.030 212.375 54.160 ;
        RECT 211.980 53.860 212.375 54.030 ;
        RECT 211.350 52.640 211.810 53.690 ;
        RECT 211.980 52.500 212.150 53.860 ;
        RECT 212.545 53.600 213.010 53.990 ;
        RECT 212.320 52.790 212.670 53.410 ;
        RECT 212.840 53.010 213.010 53.600 ;
        RECT 213.180 53.380 213.350 54.160 ;
        RECT 213.520 54.060 213.690 54.400 ;
        RECT 213.925 54.230 214.255 54.660 ;
        RECT 214.425 54.060 214.595 54.400 ;
        RECT 214.890 54.200 215.260 54.660 ;
        RECT 213.520 53.890 214.595 54.060 ;
        RECT 215.430 54.030 215.600 54.490 ;
        RECT 215.835 54.150 216.705 54.490 ;
        RECT 216.875 54.200 217.125 54.660 ;
        RECT 215.040 53.860 215.600 54.030 ;
        RECT 215.040 53.720 215.210 53.860 ;
        RECT 213.710 53.550 215.210 53.720 ;
        RECT 215.905 53.690 216.365 53.980 ;
        RECT 213.180 53.210 214.870 53.380 ;
        RECT 212.840 52.790 213.195 53.010 ;
        RECT 213.365 52.500 213.535 53.210 ;
        RECT 213.740 52.790 214.530 53.040 ;
        RECT 214.700 53.030 214.870 53.210 ;
        RECT 215.040 52.860 215.210 53.550 ;
        RECT 211.480 52.110 211.810 52.470 ;
        RECT 211.980 52.330 212.475 52.500 ;
        RECT 212.680 52.330 213.535 52.500 ;
        RECT 214.410 52.110 214.740 52.570 ;
        RECT 214.950 52.470 215.210 52.860 ;
        RECT 215.400 53.680 216.365 53.690 ;
        RECT 216.535 53.770 216.705 54.150 ;
        RECT 217.295 54.110 217.465 54.400 ;
        RECT 217.645 54.280 217.975 54.660 ;
        RECT 217.295 53.940 218.095 54.110 ;
        RECT 215.400 53.520 216.075 53.680 ;
        RECT 216.535 53.600 217.755 53.770 ;
        RECT 215.400 52.730 215.610 53.520 ;
        RECT 216.535 53.510 216.705 53.600 ;
        RECT 215.780 52.730 216.130 53.350 ;
        RECT 216.300 53.340 216.705 53.510 ;
        RECT 216.300 52.560 216.470 53.340 ;
        RECT 216.640 52.890 216.860 53.170 ;
        RECT 217.040 53.060 217.580 53.430 ;
        RECT 217.925 53.350 218.095 53.940 ;
        RECT 218.315 53.520 218.620 54.660 ;
        RECT 218.790 53.470 219.045 54.350 ;
        RECT 219.405 53.690 219.795 53.865 ;
        RECT 220.280 53.860 220.610 54.660 ;
        RECT 220.780 53.870 221.315 54.490 ;
        RECT 219.405 53.520 220.830 53.690 ;
        RECT 217.925 53.320 218.665 53.350 ;
        RECT 216.640 52.720 217.170 52.890 ;
        RECT 214.950 52.300 215.300 52.470 ;
        RECT 215.520 52.280 216.470 52.560 ;
        RECT 216.640 52.110 216.830 52.550 ;
        RECT 217.000 52.490 217.170 52.720 ;
        RECT 217.340 52.660 217.580 53.060 ;
        RECT 217.750 53.020 218.665 53.320 ;
        RECT 217.750 52.845 218.075 53.020 ;
        RECT 217.750 52.490 218.070 52.845 ;
        RECT 218.835 52.820 219.045 53.470 ;
        RECT 217.000 52.320 218.070 52.490 ;
        RECT 218.315 52.110 218.620 52.570 ;
        RECT 218.790 52.290 219.045 52.820 ;
        RECT 219.280 52.790 219.635 53.350 ;
        RECT 219.805 52.620 219.975 53.520 ;
        RECT 220.145 52.790 220.410 53.350 ;
        RECT 220.660 53.020 220.830 53.520 ;
        RECT 221.000 52.850 221.315 53.870 ;
        RECT 221.530 53.550 221.825 54.660 ;
        RECT 222.005 53.350 222.255 54.485 ;
        RECT 222.425 53.550 222.685 54.660 ;
        RECT 222.855 53.760 223.115 54.485 ;
        RECT 223.285 53.930 223.545 54.660 ;
        RECT 223.715 53.760 223.975 54.485 ;
        RECT 224.145 53.930 224.405 54.660 ;
        RECT 224.575 53.760 224.835 54.485 ;
        RECT 225.005 53.930 225.265 54.660 ;
        RECT 225.435 53.760 225.695 54.485 ;
        RECT 225.865 53.930 226.160 54.660 ;
        RECT 222.855 53.520 226.165 53.760 ;
        RECT 219.385 52.110 219.625 52.620 ;
        RECT 219.805 52.290 220.085 52.620 ;
        RECT 220.315 52.110 220.530 52.620 ;
        RECT 220.700 52.280 221.315 52.850 ;
        RECT 221.520 52.740 221.835 53.350 ;
        RECT 222.005 53.100 225.025 53.350 ;
        RECT 221.580 52.110 221.825 52.570 ;
        RECT 222.005 52.290 222.255 53.100 ;
        RECT 225.195 52.930 226.165 53.520 ;
        RECT 226.580 53.495 226.870 54.660 ;
        RECT 227.050 53.640 227.380 54.490 ;
        RECT 227.550 53.810 227.720 54.660 ;
        RECT 227.890 53.640 228.220 54.490 ;
        RECT 228.390 53.810 228.560 54.660 ;
        RECT 228.730 53.640 229.060 54.490 ;
        RECT 229.230 53.860 229.400 54.660 ;
        RECT 229.570 53.640 229.900 54.490 ;
        RECT 230.070 53.860 230.240 54.660 ;
        RECT 230.410 53.640 230.740 54.490 ;
        RECT 230.910 53.860 231.080 54.660 ;
        RECT 231.250 53.640 231.580 54.490 ;
        RECT 231.750 53.860 231.920 54.660 ;
        RECT 232.090 53.640 232.420 54.490 ;
        RECT 232.590 53.860 232.760 54.660 ;
        RECT 232.930 53.640 233.260 54.490 ;
        RECT 233.430 53.860 233.600 54.660 ;
        RECT 233.770 53.640 234.100 54.490 ;
        RECT 234.270 53.860 234.440 54.660 ;
        RECT 234.610 53.640 234.940 54.490 ;
        RECT 235.110 53.860 235.280 54.660 ;
        RECT 235.450 53.640 235.780 54.490 ;
        RECT 235.950 53.860 236.120 54.660 ;
        RECT 236.290 53.640 236.620 54.490 ;
        RECT 236.790 53.860 236.960 54.660 ;
        RECT 237.130 53.640 237.460 54.490 ;
        RECT 237.630 53.860 237.800 54.660 ;
        RECT 238.080 53.900 238.745 54.490 ;
        RECT 227.050 53.470 228.560 53.640 ;
        RECT 228.730 53.470 231.080 53.640 ;
        RECT 231.250 53.470 237.910 53.640 ;
        RECT 228.390 53.300 228.560 53.470 ;
        RECT 230.905 53.300 231.080 53.470 ;
        RECT 227.045 53.100 228.220 53.300 ;
        RECT 228.390 53.100 230.700 53.300 ;
        RECT 230.905 53.100 237.465 53.300 ;
        RECT 228.390 52.930 228.560 53.100 ;
        RECT 230.905 52.930 231.080 53.100 ;
        RECT 237.635 52.930 237.910 53.470 ;
        RECT 222.855 52.760 226.165 52.930 ;
        RECT 222.425 52.110 222.685 52.635 ;
        RECT 222.855 52.305 223.115 52.760 ;
        RECT 223.285 52.110 223.545 52.590 ;
        RECT 223.715 52.305 223.975 52.760 ;
        RECT 224.145 52.110 224.405 52.590 ;
        RECT 224.575 52.305 224.835 52.760 ;
        RECT 225.005 52.110 225.265 52.590 ;
        RECT 225.435 52.305 225.695 52.760 ;
        RECT 225.865 52.110 226.165 52.590 ;
        RECT 226.580 52.110 226.870 52.835 ;
        RECT 227.050 52.760 228.560 52.930 ;
        RECT 228.730 52.760 231.080 52.930 ;
        RECT 231.250 52.760 237.910 52.930 ;
        RECT 238.080 52.930 238.330 53.900 ;
        RECT 238.915 53.820 239.245 54.660 ;
        RECT 239.755 54.070 240.560 54.490 ;
        RECT 239.415 53.900 240.980 54.070 ;
        RECT 239.415 53.650 239.585 53.900 ;
        RECT 238.665 53.480 239.585 53.650 ;
        RECT 239.755 53.640 240.130 53.730 ;
        RECT 238.665 53.310 238.835 53.480 ;
        RECT 239.755 53.470 240.150 53.640 ;
        RECT 239.755 53.310 240.130 53.470 ;
        RECT 238.500 53.100 238.835 53.310 ;
        RECT 239.005 53.100 239.455 53.310 ;
        RECT 239.645 53.100 240.130 53.310 ;
        RECT 240.320 53.350 240.640 53.730 ;
        RECT 240.810 53.650 240.980 53.900 ;
        RECT 241.150 53.820 241.400 54.660 ;
        RECT 241.595 53.650 241.895 54.490 ;
        RECT 240.810 53.480 241.895 53.650 ;
        RECT 242.220 53.520 242.605 54.490 ;
        RECT 242.775 54.200 243.100 54.660 ;
        RECT 243.620 54.030 243.900 54.490 ;
        RECT 242.775 53.810 243.900 54.030 ;
        RECT 240.320 53.100 240.700 53.350 ;
        RECT 240.880 53.100 241.210 53.310 ;
        RECT 227.050 52.285 227.380 52.760 ;
        RECT 227.550 52.110 227.720 52.590 ;
        RECT 227.890 52.285 228.220 52.760 ;
        RECT 228.390 52.110 228.560 52.590 ;
        RECT 228.730 52.285 229.060 52.760 ;
        RECT 229.230 52.110 229.400 52.590 ;
        RECT 229.570 52.285 229.900 52.760 ;
        RECT 230.070 52.110 230.240 52.590 ;
        RECT 230.410 52.285 230.740 52.760 ;
        RECT 230.910 52.110 231.080 52.590 ;
        RECT 231.250 52.285 231.580 52.760 ;
        RECT 231.250 52.280 231.500 52.285 ;
        RECT 231.750 52.110 231.920 52.590 ;
        RECT 232.090 52.285 232.420 52.760 ;
        RECT 232.170 52.280 232.340 52.285 ;
        RECT 232.590 52.110 232.760 52.590 ;
        RECT 232.930 52.285 233.260 52.760 ;
        RECT 233.010 52.280 233.180 52.285 ;
        RECT 233.430 52.110 233.600 52.590 ;
        RECT 233.770 52.285 234.100 52.760 ;
        RECT 234.270 52.110 234.440 52.590 ;
        RECT 234.610 52.285 234.940 52.760 ;
        RECT 235.110 52.110 235.280 52.590 ;
        RECT 235.450 52.285 235.780 52.760 ;
        RECT 235.950 52.110 236.120 52.590 ;
        RECT 236.290 52.285 236.620 52.760 ;
        RECT 236.790 52.110 236.960 52.590 ;
        RECT 237.130 52.285 237.460 52.760 ;
        RECT 237.630 52.110 237.800 52.590 ;
        RECT 238.080 52.290 238.765 52.930 ;
        RECT 238.935 52.110 239.105 52.930 ;
        RECT 239.275 52.760 240.975 52.930 ;
        RECT 239.275 52.295 239.605 52.760 ;
        RECT 240.590 52.670 240.975 52.760 ;
        RECT 241.380 52.850 241.550 53.480 ;
        RECT 241.720 53.020 242.050 53.310 ;
        RECT 242.220 52.850 242.500 53.520 ;
        RECT 242.775 53.350 243.225 53.810 ;
        RECT 244.090 53.640 244.490 54.490 ;
        RECT 244.890 54.200 245.160 54.660 ;
        RECT 245.330 54.030 245.615 54.490 ;
        RECT 242.670 53.020 243.225 53.350 ;
        RECT 243.395 53.080 244.490 53.640 ;
        RECT 242.775 52.910 243.225 53.020 ;
        RECT 241.380 52.670 241.890 52.850 ;
        RECT 239.775 52.110 239.945 52.580 ;
        RECT 240.205 52.330 241.390 52.500 ;
        RECT 241.560 52.280 241.890 52.670 ;
        RECT 242.220 52.280 242.605 52.850 ;
        RECT 242.775 52.740 243.900 52.910 ;
        RECT 242.775 52.110 243.100 52.570 ;
        RECT 243.620 52.280 243.900 52.740 ;
        RECT 244.090 52.280 244.490 53.080 ;
        RECT 244.660 53.810 245.615 54.030 ;
        RECT 246.015 54.030 246.300 54.490 ;
        RECT 246.470 54.200 246.740 54.660 ;
        RECT 246.015 53.810 246.970 54.030 ;
        RECT 244.660 52.910 244.870 53.810 ;
        RECT 245.040 53.080 245.730 53.640 ;
        RECT 245.900 53.080 246.590 53.640 ;
        RECT 246.760 52.910 246.970 53.810 ;
        RECT 244.660 52.740 245.615 52.910 ;
        RECT 244.890 52.110 245.160 52.570 ;
        RECT 245.330 52.280 245.615 52.740 ;
        RECT 246.015 52.740 246.970 52.910 ;
        RECT 247.140 53.640 247.540 54.490 ;
        RECT 247.730 54.030 248.010 54.490 ;
        RECT 248.530 54.200 248.855 54.660 ;
        RECT 247.730 53.810 248.855 54.030 ;
        RECT 247.140 53.080 248.235 53.640 ;
        RECT 248.405 53.350 248.855 53.810 ;
        RECT 249.025 53.520 249.410 54.490 ;
        RECT 249.580 53.570 252.170 54.660 ;
        RECT 246.015 52.280 246.300 52.740 ;
        RECT 246.470 52.110 246.740 52.570 ;
        RECT 247.140 52.280 247.540 53.080 ;
        RECT 248.405 53.020 248.960 53.350 ;
        RECT 248.405 52.910 248.855 53.020 ;
        RECT 247.730 52.740 248.855 52.910 ;
        RECT 249.130 52.850 249.410 53.520 ;
        RECT 247.730 52.280 248.010 52.740 ;
        RECT 248.530 52.110 248.855 52.570 ;
        RECT 249.025 52.280 249.410 52.850 ;
        RECT 249.580 52.880 250.790 53.400 ;
        RECT 250.960 53.050 252.170 53.570 ;
        RECT 252.340 53.495 252.630 54.660 ;
        RECT 253.970 53.930 254.265 54.660 ;
        RECT 254.435 53.760 254.695 54.485 ;
        RECT 254.865 53.930 255.125 54.660 ;
        RECT 255.295 53.760 255.555 54.485 ;
        RECT 255.725 53.930 255.985 54.660 ;
        RECT 256.155 53.760 256.415 54.485 ;
        RECT 256.585 53.930 256.845 54.660 ;
        RECT 257.015 53.760 257.275 54.485 ;
        RECT 253.965 53.520 257.275 53.760 ;
        RECT 257.445 53.550 257.705 54.660 ;
        RECT 253.965 52.930 254.935 53.520 ;
        RECT 257.875 53.350 258.125 54.485 ;
        RECT 258.305 53.550 258.600 54.660 ;
        RECT 259.030 53.930 259.325 54.660 ;
        RECT 259.495 53.760 259.755 54.485 ;
        RECT 259.925 53.930 260.185 54.660 ;
        RECT 260.355 53.760 260.615 54.485 ;
        RECT 260.785 53.930 261.045 54.660 ;
        RECT 261.215 53.760 261.475 54.485 ;
        RECT 261.645 53.930 261.905 54.660 ;
        RECT 262.075 53.760 262.335 54.485 ;
        RECT 259.025 53.520 262.335 53.760 ;
        RECT 262.505 53.550 262.765 54.660 ;
        RECT 255.105 53.100 258.125 53.350 ;
        RECT 249.580 52.110 252.170 52.880 ;
        RECT 252.340 52.110 252.630 52.835 ;
        RECT 253.965 52.760 257.275 52.930 ;
        RECT 253.965 52.110 254.265 52.590 ;
        RECT 254.435 52.305 254.695 52.760 ;
        RECT 254.865 52.110 255.125 52.590 ;
        RECT 255.295 52.305 255.555 52.760 ;
        RECT 255.725 52.110 255.985 52.590 ;
        RECT 256.155 52.305 256.415 52.760 ;
        RECT 256.585 52.110 256.845 52.590 ;
        RECT 257.015 52.305 257.275 52.760 ;
        RECT 257.445 52.110 257.705 52.635 ;
        RECT 257.875 52.290 258.125 53.100 ;
        RECT 258.295 52.740 258.610 53.350 ;
        RECT 259.025 52.930 259.995 53.520 ;
        RECT 262.935 53.350 263.185 54.485 ;
        RECT 263.365 53.550 263.660 54.660 ;
        RECT 263.840 53.520 264.225 54.490 ;
        RECT 264.395 54.200 264.720 54.660 ;
        RECT 265.240 54.030 265.520 54.490 ;
        RECT 264.395 53.810 265.520 54.030 ;
        RECT 260.165 53.100 263.185 53.350 ;
        RECT 259.025 52.760 262.335 52.930 ;
        RECT 258.305 52.110 258.550 52.570 ;
        RECT 259.025 52.110 259.325 52.590 ;
        RECT 259.495 52.305 259.755 52.760 ;
        RECT 259.925 52.110 260.185 52.590 ;
        RECT 260.355 52.305 260.615 52.760 ;
        RECT 260.785 52.110 261.045 52.590 ;
        RECT 261.215 52.305 261.475 52.760 ;
        RECT 261.645 52.110 261.905 52.590 ;
        RECT 262.075 52.305 262.335 52.760 ;
        RECT 262.505 52.110 262.765 52.635 ;
        RECT 262.935 52.290 263.185 53.100 ;
        RECT 263.355 52.740 263.670 53.350 ;
        RECT 263.840 52.850 264.120 53.520 ;
        RECT 264.395 53.350 264.845 53.810 ;
        RECT 265.710 53.640 266.110 54.490 ;
        RECT 266.510 54.200 266.780 54.660 ;
        RECT 266.950 54.030 267.235 54.490 ;
        RECT 264.290 53.020 264.845 53.350 ;
        RECT 265.015 53.080 266.110 53.640 ;
        RECT 264.395 52.910 264.845 53.020 ;
        RECT 263.365 52.110 263.610 52.570 ;
        RECT 263.840 52.280 264.225 52.850 ;
        RECT 264.395 52.740 265.520 52.910 ;
        RECT 264.395 52.110 264.720 52.570 ;
        RECT 265.240 52.280 265.520 52.740 ;
        RECT 265.710 52.280 266.110 53.080 ;
        RECT 266.280 53.810 267.235 54.030 ;
        RECT 266.280 52.910 266.490 53.810 ;
        RECT 267.610 53.650 267.780 54.490 ;
        RECT 267.950 54.320 269.120 54.490 ;
        RECT 267.950 53.820 268.280 54.320 ;
        RECT 268.790 54.280 269.120 54.320 ;
        RECT 269.310 54.240 269.665 54.660 ;
        RECT 268.450 54.060 268.680 54.150 ;
        RECT 269.835 54.060 270.085 54.490 ;
        RECT 268.450 53.820 270.085 54.060 ;
        RECT 270.255 53.900 270.585 54.660 ;
        RECT 270.755 53.820 271.010 54.490 ;
        RECT 266.660 53.080 267.350 53.640 ;
        RECT 267.610 53.480 270.670 53.650 ;
        RECT 267.525 53.100 267.875 53.310 ;
        RECT 268.045 53.100 268.490 53.300 ;
        RECT 268.660 53.100 269.135 53.300 ;
        RECT 266.280 52.740 267.235 52.910 ;
        RECT 266.510 52.110 266.780 52.570 ;
        RECT 266.950 52.280 267.235 52.740 ;
        RECT 267.610 52.760 268.675 52.930 ;
        RECT 267.610 52.280 267.780 52.760 ;
        RECT 267.950 52.110 268.280 52.590 ;
        RECT 268.505 52.530 268.675 52.760 ;
        RECT 268.855 52.700 269.135 53.100 ;
        RECT 269.405 53.100 269.735 53.300 ;
        RECT 269.905 53.100 270.270 53.300 ;
        RECT 269.405 52.700 269.690 53.100 ;
        RECT 270.500 52.930 270.670 53.480 ;
        RECT 269.870 52.760 270.670 52.930 ;
        RECT 269.870 52.530 270.040 52.760 ;
        RECT 270.840 52.690 271.010 53.820 ;
        RECT 271.200 53.570 274.710 54.660 ;
        RECT 270.825 52.620 271.010 52.690 ;
        RECT 270.800 52.610 271.010 52.620 ;
        RECT 268.505 52.280 270.040 52.530 ;
        RECT 270.210 52.110 270.540 52.590 ;
        RECT 270.755 52.280 271.010 52.610 ;
        RECT 271.200 52.880 272.850 53.400 ;
        RECT 273.020 53.050 274.710 53.570 ;
        RECT 274.925 53.520 275.220 54.660 ;
        RECT 275.480 53.690 275.810 54.490 ;
        RECT 275.980 53.860 276.150 54.660 ;
        RECT 276.320 53.690 276.650 54.490 ;
        RECT 276.820 53.860 276.990 54.660 ;
        RECT 277.160 53.710 277.490 54.490 ;
        RECT 277.660 54.200 277.830 54.660 ;
        RECT 277.160 53.690 277.930 53.710 ;
        RECT 275.480 53.520 277.930 53.690 ;
        RECT 274.900 53.100 277.410 53.350 ;
        RECT 277.580 52.930 277.930 53.520 ;
        RECT 278.100 53.495 278.390 54.660 ;
        RECT 271.200 52.110 274.710 52.880 ;
        RECT 275.560 52.750 277.930 52.930 ;
        RECT 278.565 53.470 278.820 54.350 ;
        RECT 278.990 53.520 279.295 54.660 ;
        RECT 279.635 54.280 279.965 54.660 ;
        RECT 280.145 54.110 280.315 54.400 ;
        RECT 280.485 54.200 280.735 54.660 ;
        RECT 279.515 53.940 280.315 54.110 ;
        RECT 280.905 54.150 281.775 54.490 ;
        RECT 274.925 52.110 275.190 52.570 ;
        RECT 275.560 52.280 275.730 52.750 ;
        RECT 275.980 52.110 276.150 52.570 ;
        RECT 276.400 52.280 276.570 52.750 ;
        RECT 276.820 52.110 276.990 52.570 ;
        RECT 277.240 52.280 277.410 52.750 ;
        RECT 277.580 52.110 277.830 52.575 ;
        RECT 278.100 52.110 278.390 52.835 ;
        RECT 278.565 52.820 278.775 53.470 ;
        RECT 279.515 53.350 279.685 53.940 ;
        RECT 280.905 53.770 281.075 54.150 ;
        RECT 282.010 54.030 282.180 54.490 ;
        RECT 282.350 54.200 282.720 54.660 ;
        RECT 283.015 54.060 283.185 54.400 ;
        RECT 283.355 54.230 283.685 54.660 ;
        RECT 283.920 54.060 284.090 54.400 ;
        RECT 279.855 53.600 281.075 53.770 ;
        RECT 281.245 53.690 281.705 53.980 ;
        RECT 282.010 53.860 282.570 54.030 ;
        RECT 283.015 53.890 284.090 54.060 ;
        RECT 284.260 54.160 284.940 54.490 ;
        RECT 285.155 54.160 285.405 54.490 ;
        RECT 285.575 54.200 285.825 54.660 ;
        RECT 282.400 53.720 282.570 53.860 ;
        RECT 281.245 53.680 282.210 53.690 ;
        RECT 280.905 53.510 281.075 53.600 ;
        RECT 281.535 53.520 282.210 53.680 ;
        RECT 278.945 53.320 279.685 53.350 ;
        RECT 278.945 53.020 279.860 53.320 ;
        RECT 279.535 52.845 279.860 53.020 ;
        RECT 278.565 52.290 278.820 52.820 ;
        RECT 278.990 52.110 279.295 52.570 ;
        RECT 279.540 52.490 279.860 52.845 ;
        RECT 280.030 53.060 280.570 53.430 ;
        RECT 280.905 53.340 281.310 53.510 ;
        RECT 280.030 52.660 280.270 53.060 ;
        RECT 280.750 52.890 280.970 53.170 ;
        RECT 280.440 52.720 280.970 52.890 ;
        RECT 280.440 52.490 280.610 52.720 ;
        RECT 281.140 52.560 281.310 53.340 ;
        RECT 281.480 52.730 281.830 53.350 ;
        RECT 282.000 52.730 282.210 53.520 ;
        RECT 282.400 53.550 283.900 53.720 ;
        RECT 282.400 52.860 282.570 53.550 ;
        RECT 284.260 53.380 284.430 54.160 ;
        RECT 285.235 54.030 285.405 54.160 ;
        RECT 282.740 53.210 284.430 53.380 ;
        RECT 284.600 53.600 285.065 53.990 ;
        RECT 285.235 53.860 285.630 54.030 ;
        RECT 282.740 53.030 282.910 53.210 ;
        RECT 279.540 52.320 280.610 52.490 ;
        RECT 280.780 52.110 280.970 52.550 ;
        RECT 281.140 52.280 282.090 52.560 ;
        RECT 282.400 52.470 282.660 52.860 ;
        RECT 283.080 52.790 283.870 53.040 ;
        RECT 282.310 52.300 282.660 52.470 ;
        RECT 282.870 52.110 283.200 52.570 ;
        RECT 284.075 52.500 284.245 53.210 ;
        RECT 284.600 53.010 284.770 53.600 ;
        RECT 284.415 52.790 284.770 53.010 ;
        RECT 284.940 52.790 285.290 53.410 ;
        RECT 285.460 52.500 285.630 53.860 ;
        RECT 285.995 53.690 286.320 54.475 ;
        RECT 285.800 52.640 286.260 53.690 ;
        RECT 284.075 52.330 284.930 52.500 ;
        RECT 285.135 52.330 285.630 52.500 ;
        RECT 285.800 52.110 286.130 52.470 ;
        RECT 286.490 52.370 286.660 54.490 ;
        RECT 286.830 54.160 287.160 54.660 ;
        RECT 287.330 53.990 287.585 54.490 ;
        RECT 286.835 53.820 287.585 53.990 ;
        RECT 286.835 52.830 287.065 53.820 ;
        RECT 287.235 53.000 287.585 53.650 ;
        RECT 287.770 53.550 288.065 54.660 ;
        RECT 288.245 53.350 288.495 54.485 ;
        RECT 288.665 53.550 288.925 54.660 ;
        RECT 289.095 53.760 289.355 54.485 ;
        RECT 289.525 53.930 289.785 54.660 ;
        RECT 289.955 53.760 290.215 54.485 ;
        RECT 290.385 53.930 290.645 54.660 ;
        RECT 290.815 53.760 291.075 54.485 ;
        RECT 291.245 53.930 291.505 54.660 ;
        RECT 291.675 53.760 291.935 54.485 ;
        RECT 292.105 53.930 292.400 54.660 ;
        RECT 292.820 54.225 298.165 54.660 ;
        RECT 289.095 53.520 292.405 53.760 ;
        RECT 286.835 52.660 287.585 52.830 ;
        RECT 287.760 52.740 288.075 53.350 ;
        RECT 288.245 53.100 291.265 53.350 ;
        RECT 286.830 52.110 287.160 52.490 ;
        RECT 287.330 52.370 287.585 52.660 ;
        RECT 287.820 52.110 288.065 52.570 ;
        RECT 288.245 52.290 288.495 53.100 ;
        RECT 291.435 52.930 292.405 53.520 ;
        RECT 289.095 52.760 292.405 52.930 ;
        RECT 288.665 52.110 288.925 52.635 ;
        RECT 289.095 52.305 289.355 52.760 ;
        RECT 289.525 52.110 289.785 52.590 ;
        RECT 289.955 52.305 290.215 52.760 ;
        RECT 290.385 52.110 290.645 52.590 ;
        RECT 290.815 52.305 291.075 52.760 ;
        RECT 291.245 52.110 291.505 52.590 ;
        RECT 291.675 52.305 291.935 52.760 ;
        RECT 294.405 52.655 294.745 53.485 ;
        RECT 296.225 52.975 296.575 54.225 ;
        RECT 298.340 53.570 300.930 54.660 ;
        RECT 298.340 52.880 299.550 53.400 ;
        RECT 299.720 53.050 300.930 53.570 ;
        RECT 301.100 53.690 301.410 54.490 ;
        RECT 301.580 53.860 301.890 54.660 ;
        RECT 302.060 54.030 302.320 54.490 ;
        RECT 302.490 54.200 302.745 54.660 ;
        RECT 302.920 54.030 303.180 54.490 ;
        RECT 302.060 53.860 303.180 54.030 ;
        RECT 301.100 53.520 302.130 53.690 ;
        RECT 292.105 52.110 292.405 52.590 ;
        RECT 292.820 52.110 298.165 52.655 ;
        RECT 298.340 52.110 300.930 52.880 ;
        RECT 301.100 52.610 301.270 53.520 ;
        RECT 301.440 52.780 301.790 53.350 ;
        RECT 301.960 53.270 302.130 53.520 ;
        RECT 302.920 53.610 303.180 53.860 ;
        RECT 303.350 53.790 303.635 54.660 ;
        RECT 302.920 53.440 303.675 53.610 ;
        RECT 303.860 53.495 304.150 54.660 ;
        RECT 304.435 54.030 304.720 54.490 ;
        RECT 304.890 54.200 305.160 54.660 ;
        RECT 304.435 53.810 305.390 54.030 ;
        RECT 301.960 53.100 303.100 53.270 ;
        RECT 303.270 52.930 303.675 53.440 ;
        RECT 304.320 53.080 305.010 53.640 ;
        RECT 302.025 52.760 303.675 52.930 ;
        RECT 305.180 52.910 305.390 53.810 ;
        RECT 301.100 52.280 301.400 52.610 ;
        RECT 301.570 52.110 301.845 52.590 ;
        RECT 302.025 52.370 302.320 52.760 ;
        RECT 302.490 52.110 302.745 52.590 ;
        RECT 302.920 52.370 303.180 52.760 ;
        RECT 303.350 52.110 303.630 52.590 ;
        RECT 303.860 52.110 304.150 52.835 ;
        RECT 304.435 52.740 305.390 52.910 ;
        RECT 305.560 53.640 305.960 54.490 ;
        RECT 306.150 54.030 306.430 54.490 ;
        RECT 306.950 54.200 307.275 54.660 ;
        RECT 306.150 53.810 307.275 54.030 ;
        RECT 305.560 53.080 306.655 53.640 ;
        RECT 306.825 53.350 307.275 53.810 ;
        RECT 307.445 53.520 307.830 54.490 ;
        RECT 304.435 52.280 304.720 52.740 ;
        RECT 304.890 52.110 305.160 52.570 ;
        RECT 305.560 52.280 305.960 53.080 ;
        RECT 306.825 53.020 307.380 53.350 ;
        RECT 306.825 52.910 307.275 53.020 ;
        RECT 306.150 52.740 307.275 52.910 ;
        RECT 307.550 52.850 307.830 53.520 ;
        RECT 306.150 52.280 306.430 52.740 ;
        RECT 306.950 52.110 307.275 52.570 ;
        RECT 307.445 52.280 307.830 52.850 ;
        RECT 308.460 53.585 308.730 54.490 ;
        RECT 308.900 53.900 309.230 54.660 ;
        RECT 309.410 53.730 309.580 54.490 ;
        RECT 308.460 52.785 308.630 53.585 ;
        RECT 308.915 53.560 309.580 53.730 ;
        RECT 309.840 53.570 311.050 54.660 ;
        RECT 308.915 53.415 309.085 53.560 ;
        RECT 308.800 53.085 309.085 53.415 ;
        RECT 308.915 52.830 309.085 53.085 ;
        RECT 309.320 53.010 309.650 53.380 ;
        RECT 309.840 53.030 310.360 53.570 ;
        RECT 310.530 52.860 311.050 53.400 ;
        RECT 308.460 52.280 308.720 52.785 ;
        RECT 308.915 52.660 309.580 52.830 ;
        RECT 308.900 52.110 309.230 52.490 ;
        RECT 309.410 52.280 309.580 52.660 ;
        RECT 309.840 52.110 311.050 52.860 ;
        RECT 162.095 51.940 311.135 52.110 ;
        RECT 162.180 51.190 163.390 51.940 ;
        RECT 162.180 50.650 162.700 51.190 ;
        RECT 163.560 51.170 165.230 51.940 ;
        RECT 165.865 51.390 166.120 51.680 ;
        RECT 166.290 51.560 166.620 51.940 ;
        RECT 165.865 51.220 166.615 51.390 ;
        RECT 162.870 50.480 163.390 51.020 ;
        RECT 163.560 50.650 164.310 51.170 ;
        RECT 164.480 50.480 165.230 51.000 ;
        RECT 162.180 49.390 163.390 50.480 ;
        RECT 163.560 49.390 165.230 50.480 ;
        RECT 165.865 50.400 166.215 51.050 ;
        RECT 166.385 50.230 166.615 51.220 ;
        RECT 165.865 50.060 166.615 50.230 ;
        RECT 165.865 49.560 166.120 50.060 ;
        RECT 166.290 49.390 166.620 49.890 ;
        RECT 166.790 49.560 166.960 51.680 ;
        RECT 167.320 51.580 167.650 51.940 ;
        RECT 167.820 51.550 168.315 51.720 ;
        RECT 168.520 51.550 169.375 51.720 ;
        RECT 167.190 50.360 167.650 51.410 ;
        RECT 167.130 49.575 167.455 50.360 ;
        RECT 167.820 50.190 167.990 51.550 ;
        RECT 168.160 50.640 168.510 51.260 ;
        RECT 168.680 51.040 169.035 51.260 ;
        RECT 168.680 50.450 168.850 51.040 ;
        RECT 169.205 50.840 169.375 51.550 ;
        RECT 170.250 51.480 170.580 51.940 ;
        RECT 170.790 51.580 171.140 51.750 ;
        RECT 169.580 51.010 170.370 51.260 ;
        RECT 170.790 51.190 171.050 51.580 ;
        RECT 171.360 51.490 172.310 51.770 ;
        RECT 172.480 51.500 172.670 51.940 ;
        RECT 172.840 51.560 173.910 51.730 ;
        RECT 170.540 50.840 170.710 51.020 ;
        RECT 167.820 50.020 168.215 50.190 ;
        RECT 168.385 50.060 168.850 50.450 ;
        RECT 169.020 50.670 170.710 50.840 ;
        RECT 168.045 49.890 168.215 50.020 ;
        RECT 169.020 49.890 169.190 50.670 ;
        RECT 170.880 50.500 171.050 51.190 ;
        RECT 169.550 50.330 171.050 50.500 ;
        RECT 171.240 50.530 171.450 51.320 ;
        RECT 171.620 50.700 171.970 51.320 ;
        RECT 172.140 50.710 172.310 51.490 ;
        RECT 172.840 51.330 173.010 51.560 ;
        RECT 172.480 51.160 173.010 51.330 ;
        RECT 172.480 50.880 172.700 51.160 ;
        RECT 173.180 50.990 173.420 51.390 ;
        RECT 172.140 50.540 172.545 50.710 ;
        RECT 172.880 50.620 173.420 50.990 ;
        RECT 173.590 51.205 173.910 51.560 ;
        RECT 174.155 51.480 174.460 51.940 ;
        RECT 174.630 51.230 174.885 51.760 ;
        RECT 173.590 51.030 173.915 51.205 ;
        RECT 173.590 50.730 174.505 51.030 ;
        RECT 173.765 50.700 174.505 50.730 ;
        RECT 171.240 50.370 171.915 50.530 ;
        RECT 172.375 50.450 172.545 50.540 ;
        RECT 171.240 50.360 172.205 50.370 ;
        RECT 170.880 50.190 171.050 50.330 ;
        RECT 167.625 49.390 167.875 49.850 ;
        RECT 168.045 49.560 168.295 49.890 ;
        RECT 168.510 49.560 169.190 49.890 ;
        RECT 169.360 49.990 170.435 50.160 ;
        RECT 170.880 50.020 171.440 50.190 ;
        RECT 171.745 50.070 172.205 50.360 ;
        RECT 172.375 50.280 173.595 50.450 ;
        RECT 169.360 49.650 169.530 49.990 ;
        RECT 169.765 49.390 170.095 49.820 ;
        RECT 170.265 49.650 170.435 49.990 ;
        RECT 170.730 49.390 171.100 49.850 ;
        RECT 171.270 49.560 171.440 50.020 ;
        RECT 172.375 49.900 172.545 50.280 ;
        RECT 173.765 50.110 173.935 50.700 ;
        RECT 174.675 50.580 174.885 51.230 ;
        RECT 175.065 51.390 175.320 51.680 ;
        RECT 175.490 51.560 175.820 51.940 ;
        RECT 175.065 51.220 175.815 51.390 ;
        RECT 171.675 49.560 172.545 49.900 ;
        RECT 173.135 49.940 173.935 50.110 ;
        RECT 172.715 49.390 172.965 49.850 ;
        RECT 173.135 49.650 173.305 49.940 ;
        RECT 173.485 49.390 173.815 49.770 ;
        RECT 174.155 49.390 174.460 50.530 ;
        RECT 174.630 49.700 174.885 50.580 ;
        RECT 175.065 50.400 175.415 51.050 ;
        RECT 175.585 50.230 175.815 51.220 ;
        RECT 175.065 50.060 175.815 50.230 ;
        RECT 175.065 49.560 175.320 50.060 ;
        RECT 175.490 49.390 175.820 49.890 ;
        RECT 175.990 49.560 176.160 51.680 ;
        RECT 176.520 51.580 176.850 51.940 ;
        RECT 177.020 51.550 177.515 51.720 ;
        RECT 177.720 51.550 178.575 51.720 ;
        RECT 176.390 50.360 176.850 51.410 ;
        RECT 176.330 49.575 176.655 50.360 ;
        RECT 177.020 50.190 177.190 51.550 ;
        RECT 177.360 50.640 177.710 51.260 ;
        RECT 177.880 51.040 178.235 51.260 ;
        RECT 177.880 50.450 178.050 51.040 ;
        RECT 178.405 50.840 178.575 51.550 ;
        RECT 179.450 51.480 179.780 51.940 ;
        RECT 179.990 51.580 180.340 51.750 ;
        RECT 178.780 51.010 179.570 51.260 ;
        RECT 179.990 51.190 180.250 51.580 ;
        RECT 180.560 51.490 181.510 51.770 ;
        RECT 181.680 51.500 181.870 51.940 ;
        RECT 182.040 51.560 183.110 51.730 ;
        RECT 179.740 50.840 179.910 51.020 ;
        RECT 177.020 50.020 177.415 50.190 ;
        RECT 177.585 50.060 178.050 50.450 ;
        RECT 178.220 50.670 179.910 50.840 ;
        RECT 177.245 49.890 177.415 50.020 ;
        RECT 178.220 49.890 178.390 50.670 ;
        RECT 180.080 50.500 180.250 51.190 ;
        RECT 178.750 50.330 180.250 50.500 ;
        RECT 180.440 50.530 180.650 51.320 ;
        RECT 180.820 50.700 181.170 51.320 ;
        RECT 181.340 50.710 181.510 51.490 ;
        RECT 182.040 51.330 182.210 51.560 ;
        RECT 181.680 51.160 182.210 51.330 ;
        RECT 181.680 50.880 181.900 51.160 ;
        RECT 182.380 50.990 182.620 51.390 ;
        RECT 181.340 50.540 181.745 50.710 ;
        RECT 182.080 50.620 182.620 50.990 ;
        RECT 182.790 51.205 183.110 51.560 ;
        RECT 183.355 51.480 183.660 51.940 ;
        RECT 183.830 51.230 184.085 51.760 ;
        RECT 184.265 51.685 184.600 51.730 ;
        RECT 182.790 51.030 183.115 51.205 ;
        RECT 182.790 50.730 183.705 51.030 ;
        RECT 182.965 50.700 183.705 50.730 ;
        RECT 180.440 50.370 181.115 50.530 ;
        RECT 181.575 50.450 181.745 50.540 ;
        RECT 180.440 50.360 181.405 50.370 ;
        RECT 180.080 50.190 180.250 50.330 ;
        RECT 176.825 49.390 177.075 49.850 ;
        RECT 177.245 49.560 177.495 49.890 ;
        RECT 177.710 49.560 178.390 49.890 ;
        RECT 178.560 49.990 179.635 50.160 ;
        RECT 180.080 50.020 180.640 50.190 ;
        RECT 180.945 50.070 181.405 50.360 ;
        RECT 181.575 50.280 182.795 50.450 ;
        RECT 178.560 49.650 178.730 49.990 ;
        RECT 178.965 49.390 179.295 49.820 ;
        RECT 179.465 49.650 179.635 49.990 ;
        RECT 179.930 49.390 180.300 49.850 ;
        RECT 180.470 49.560 180.640 50.020 ;
        RECT 181.575 49.900 181.745 50.280 ;
        RECT 182.965 50.110 183.135 50.700 ;
        RECT 183.875 50.580 184.085 51.230 ;
        RECT 180.875 49.560 181.745 49.900 ;
        RECT 182.335 49.940 183.135 50.110 ;
        RECT 181.915 49.390 182.165 49.850 ;
        RECT 182.335 49.650 182.505 49.940 ;
        RECT 182.685 49.390 183.015 49.770 ;
        RECT 183.355 49.390 183.660 50.530 ;
        RECT 183.830 49.700 184.085 50.580 ;
        RECT 184.260 51.220 184.600 51.685 ;
        RECT 184.770 51.560 185.100 51.940 ;
        RECT 184.260 50.530 184.430 51.220 ;
        RECT 184.600 50.700 184.860 51.030 ;
        RECT 184.260 49.560 184.520 50.530 ;
        RECT 184.690 50.150 184.860 50.700 ;
        RECT 185.030 50.330 185.370 51.360 ;
        RECT 185.560 50.580 185.830 51.605 ;
        RECT 185.560 50.410 185.870 50.580 ;
        RECT 185.560 50.330 185.830 50.410 ;
        RECT 186.055 50.330 186.335 51.605 ;
        RECT 186.535 51.440 186.765 51.770 ;
        RECT 187.010 51.560 187.340 51.940 ;
        RECT 186.535 50.150 186.705 51.440 ;
        RECT 187.510 51.370 187.685 51.770 ;
        RECT 187.055 51.200 187.685 51.370 ;
        RECT 187.940 51.215 188.230 51.940 ;
        RECT 189.405 51.440 189.900 51.770 ;
        RECT 187.055 51.030 187.225 51.200 ;
        RECT 186.875 50.700 187.225 51.030 ;
        RECT 184.690 49.980 186.705 50.150 ;
        RECT 187.055 50.180 187.225 50.700 ;
        RECT 187.405 50.350 187.770 51.030 ;
        RECT 187.055 50.010 187.685 50.180 ;
        RECT 184.715 49.390 185.045 49.800 ;
        RECT 185.245 49.560 185.415 49.980 ;
        RECT 185.630 49.390 186.300 49.800 ;
        RECT 186.535 49.560 186.705 49.980 ;
        RECT 187.010 49.390 187.340 49.830 ;
        RECT 187.510 49.560 187.685 50.010 ;
        RECT 187.940 49.390 188.230 50.555 ;
        RECT 189.320 49.950 189.560 51.260 ;
        RECT 189.730 50.530 189.900 51.440 ;
        RECT 190.120 50.700 190.470 51.665 ;
        RECT 190.650 50.700 190.950 51.670 ;
        RECT 191.130 50.700 191.410 51.670 ;
        RECT 191.590 51.140 191.860 51.940 ;
        RECT 192.030 51.220 192.370 51.730 ;
        RECT 193.935 51.415 194.230 51.940 ;
        RECT 191.605 50.700 191.935 50.950 ;
        RECT 191.605 50.530 191.920 50.700 ;
        RECT 189.730 50.360 191.920 50.530 ;
        RECT 189.325 49.390 189.660 49.770 ;
        RECT 189.830 49.560 190.080 50.360 ;
        RECT 190.300 49.390 190.630 50.110 ;
        RECT 190.815 49.560 191.065 50.360 ;
        RECT 191.530 49.390 191.860 50.190 ;
        RECT 192.110 49.820 192.370 51.220 ;
        RECT 194.400 51.300 194.625 51.745 ;
        RECT 194.795 51.470 195.125 51.940 ;
        RECT 195.305 51.390 195.560 51.680 ;
        RECT 195.730 51.560 196.060 51.940 ;
        RECT 194.400 51.130 195.130 51.300 ;
        RECT 195.305 51.220 196.055 51.390 ;
        RECT 193.460 50.735 194.680 50.960 ;
        RECT 194.850 50.565 195.130 51.130 ;
        RECT 192.030 49.560 192.370 49.820 ;
        RECT 193.530 50.395 195.130 50.565 ;
        RECT 195.305 50.400 195.655 51.050 ;
        RECT 193.530 49.590 193.785 50.395 ;
        RECT 193.955 49.390 194.215 50.225 ;
        RECT 194.385 49.590 194.645 50.395 ;
        RECT 195.825 50.230 196.055 51.220 ;
        RECT 194.815 49.390 195.070 50.225 ;
        RECT 195.305 50.060 196.055 50.230 ;
        RECT 195.305 49.560 195.560 50.060 ;
        RECT 195.730 49.390 196.060 49.890 ;
        RECT 196.230 49.560 196.400 51.680 ;
        RECT 196.760 51.580 197.090 51.940 ;
        RECT 197.260 51.550 197.755 51.720 ;
        RECT 197.960 51.550 198.815 51.720 ;
        RECT 196.630 50.360 197.090 51.410 ;
        RECT 196.570 49.575 196.895 50.360 ;
        RECT 197.260 50.190 197.430 51.550 ;
        RECT 197.600 50.640 197.950 51.260 ;
        RECT 198.120 51.040 198.475 51.260 ;
        RECT 198.120 50.450 198.290 51.040 ;
        RECT 198.645 50.840 198.815 51.550 ;
        RECT 199.690 51.480 200.020 51.940 ;
        RECT 200.230 51.580 200.580 51.750 ;
        RECT 199.020 51.010 199.810 51.260 ;
        RECT 200.230 51.190 200.490 51.580 ;
        RECT 200.800 51.490 201.750 51.770 ;
        RECT 201.920 51.500 202.110 51.940 ;
        RECT 202.280 51.560 203.350 51.730 ;
        RECT 199.980 50.840 200.150 51.020 ;
        RECT 197.260 50.020 197.655 50.190 ;
        RECT 197.825 50.060 198.290 50.450 ;
        RECT 198.460 50.670 200.150 50.840 ;
        RECT 197.485 49.890 197.655 50.020 ;
        RECT 198.460 49.890 198.630 50.670 ;
        RECT 200.320 50.500 200.490 51.190 ;
        RECT 198.990 50.330 200.490 50.500 ;
        RECT 200.680 50.530 200.890 51.320 ;
        RECT 201.060 50.700 201.410 51.320 ;
        RECT 201.580 50.710 201.750 51.490 ;
        RECT 202.280 51.330 202.450 51.560 ;
        RECT 201.920 51.160 202.450 51.330 ;
        RECT 201.920 50.880 202.140 51.160 ;
        RECT 202.620 50.990 202.860 51.390 ;
        RECT 201.580 50.540 201.985 50.710 ;
        RECT 202.320 50.620 202.860 50.990 ;
        RECT 203.030 51.205 203.350 51.560 ;
        RECT 203.595 51.480 203.900 51.940 ;
        RECT 204.070 51.230 204.325 51.760 ;
        RECT 203.030 51.030 203.355 51.205 ;
        RECT 203.030 50.730 203.945 51.030 ;
        RECT 203.205 50.700 203.945 50.730 ;
        RECT 200.680 50.370 201.355 50.530 ;
        RECT 201.815 50.450 201.985 50.540 ;
        RECT 200.680 50.360 201.645 50.370 ;
        RECT 200.320 50.190 200.490 50.330 ;
        RECT 197.065 49.390 197.315 49.850 ;
        RECT 197.485 49.560 197.735 49.890 ;
        RECT 197.950 49.560 198.630 49.890 ;
        RECT 198.800 49.990 199.875 50.160 ;
        RECT 200.320 50.020 200.880 50.190 ;
        RECT 201.185 50.070 201.645 50.360 ;
        RECT 201.815 50.280 203.035 50.450 ;
        RECT 198.800 49.650 198.970 49.990 ;
        RECT 199.205 49.390 199.535 49.820 ;
        RECT 199.705 49.650 199.875 49.990 ;
        RECT 200.170 49.390 200.540 49.850 ;
        RECT 200.710 49.560 200.880 50.020 ;
        RECT 201.815 49.900 201.985 50.280 ;
        RECT 203.205 50.110 203.375 50.700 ;
        RECT 204.115 50.580 204.325 51.230 ;
        RECT 204.505 51.390 204.760 51.680 ;
        RECT 204.930 51.560 205.260 51.940 ;
        RECT 204.505 51.220 205.255 51.390 ;
        RECT 201.115 49.560 201.985 49.900 ;
        RECT 202.575 49.940 203.375 50.110 ;
        RECT 202.155 49.390 202.405 49.850 ;
        RECT 202.575 49.650 202.745 49.940 ;
        RECT 202.925 49.390 203.255 49.770 ;
        RECT 203.595 49.390 203.900 50.530 ;
        RECT 204.070 49.700 204.325 50.580 ;
        RECT 204.505 50.400 204.855 51.050 ;
        RECT 205.025 50.230 205.255 51.220 ;
        RECT 204.505 50.060 205.255 50.230 ;
        RECT 204.505 49.560 204.760 50.060 ;
        RECT 204.930 49.390 205.260 49.890 ;
        RECT 205.430 49.560 205.600 51.680 ;
        RECT 205.960 51.580 206.290 51.940 ;
        RECT 206.460 51.550 206.955 51.720 ;
        RECT 207.160 51.550 208.015 51.720 ;
        RECT 205.830 50.360 206.290 51.410 ;
        RECT 205.770 49.575 206.095 50.360 ;
        RECT 206.460 50.190 206.630 51.550 ;
        RECT 206.800 50.640 207.150 51.260 ;
        RECT 207.320 51.040 207.675 51.260 ;
        RECT 207.320 50.450 207.490 51.040 ;
        RECT 207.845 50.840 208.015 51.550 ;
        RECT 208.890 51.480 209.220 51.940 ;
        RECT 209.430 51.580 209.780 51.750 ;
        RECT 208.220 51.010 209.010 51.260 ;
        RECT 209.430 51.190 209.690 51.580 ;
        RECT 210.000 51.490 210.950 51.770 ;
        RECT 211.120 51.500 211.310 51.940 ;
        RECT 211.480 51.560 212.550 51.730 ;
        RECT 209.180 50.840 209.350 51.020 ;
        RECT 206.460 50.020 206.855 50.190 ;
        RECT 207.025 50.060 207.490 50.450 ;
        RECT 207.660 50.670 209.350 50.840 ;
        RECT 206.685 49.890 206.855 50.020 ;
        RECT 207.660 49.890 207.830 50.670 ;
        RECT 209.520 50.500 209.690 51.190 ;
        RECT 208.190 50.330 209.690 50.500 ;
        RECT 209.880 50.530 210.090 51.320 ;
        RECT 210.260 50.700 210.610 51.320 ;
        RECT 210.780 50.710 210.950 51.490 ;
        RECT 211.480 51.330 211.650 51.560 ;
        RECT 211.120 51.160 211.650 51.330 ;
        RECT 211.120 50.880 211.340 51.160 ;
        RECT 211.820 50.990 212.060 51.390 ;
        RECT 210.780 50.540 211.185 50.710 ;
        RECT 211.520 50.620 212.060 50.990 ;
        RECT 212.230 51.205 212.550 51.560 ;
        RECT 212.795 51.480 213.100 51.940 ;
        RECT 213.270 51.230 213.525 51.760 ;
        RECT 212.230 51.030 212.555 51.205 ;
        RECT 212.230 50.730 213.145 51.030 ;
        RECT 212.405 50.700 213.145 50.730 ;
        RECT 209.880 50.370 210.555 50.530 ;
        RECT 211.015 50.450 211.185 50.540 ;
        RECT 209.880 50.360 210.845 50.370 ;
        RECT 209.520 50.190 209.690 50.330 ;
        RECT 206.265 49.390 206.515 49.850 ;
        RECT 206.685 49.560 206.935 49.890 ;
        RECT 207.150 49.560 207.830 49.890 ;
        RECT 208.000 49.990 209.075 50.160 ;
        RECT 209.520 50.020 210.080 50.190 ;
        RECT 210.385 50.070 210.845 50.360 ;
        RECT 211.015 50.280 212.235 50.450 ;
        RECT 208.000 49.650 208.170 49.990 ;
        RECT 208.405 49.390 208.735 49.820 ;
        RECT 208.905 49.650 209.075 49.990 ;
        RECT 209.370 49.390 209.740 49.850 ;
        RECT 209.910 49.560 210.080 50.020 ;
        RECT 211.015 49.900 211.185 50.280 ;
        RECT 212.405 50.110 212.575 50.700 ;
        RECT 213.315 50.580 213.525 51.230 ;
        RECT 213.700 51.215 213.990 51.940 ;
        RECT 214.165 51.390 214.420 51.680 ;
        RECT 214.590 51.560 214.920 51.940 ;
        RECT 214.165 51.220 214.915 51.390 ;
        RECT 210.315 49.560 211.185 49.900 ;
        RECT 211.775 49.940 212.575 50.110 ;
        RECT 211.355 49.390 211.605 49.850 ;
        RECT 211.775 49.650 211.945 49.940 ;
        RECT 212.125 49.390 212.455 49.770 ;
        RECT 212.795 49.390 213.100 50.530 ;
        RECT 213.270 49.700 213.525 50.580 ;
        RECT 213.700 49.390 213.990 50.555 ;
        RECT 214.165 50.400 214.515 51.050 ;
        RECT 214.685 50.230 214.915 51.220 ;
        RECT 214.165 50.060 214.915 50.230 ;
        RECT 214.165 49.560 214.420 50.060 ;
        RECT 214.590 49.390 214.920 49.890 ;
        RECT 215.090 49.560 215.260 51.680 ;
        RECT 215.620 51.580 215.950 51.940 ;
        RECT 216.120 51.550 216.615 51.720 ;
        RECT 216.820 51.550 217.675 51.720 ;
        RECT 215.490 50.360 215.950 51.410 ;
        RECT 215.430 49.575 215.755 50.360 ;
        RECT 216.120 50.190 216.290 51.550 ;
        RECT 216.460 50.640 216.810 51.260 ;
        RECT 216.980 51.040 217.335 51.260 ;
        RECT 216.980 50.450 217.150 51.040 ;
        RECT 217.505 50.840 217.675 51.550 ;
        RECT 218.550 51.480 218.880 51.940 ;
        RECT 219.090 51.580 219.440 51.750 ;
        RECT 217.880 51.010 218.670 51.260 ;
        RECT 219.090 51.190 219.350 51.580 ;
        RECT 219.660 51.490 220.610 51.770 ;
        RECT 220.780 51.500 220.970 51.940 ;
        RECT 221.140 51.560 222.210 51.730 ;
        RECT 218.840 50.840 219.010 51.020 ;
        RECT 216.120 50.020 216.515 50.190 ;
        RECT 216.685 50.060 217.150 50.450 ;
        RECT 217.320 50.670 219.010 50.840 ;
        RECT 216.345 49.890 216.515 50.020 ;
        RECT 217.320 49.890 217.490 50.670 ;
        RECT 219.180 50.500 219.350 51.190 ;
        RECT 217.850 50.330 219.350 50.500 ;
        RECT 219.540 50.530 219.750 51.320 ;
        RECT 219.920 50.700 220.270 51.320 ;
        RECT 220.440 50.710 220.610 51.490 ;
        RECT 221.140 51.330 221.310 51.560 ;
        RECT 220.780 51.160 221.310 51.330 ;
        RECT 220.780 50.880 221.000 51.160 ;
        RECT 221.480 50.990 221.720 51.390 ;
        RECT 220.440 50.540 220.845 50.710 ;
        RECT 221.180 50.620 221.720 50.990 ;
        RECT 221.890 51.205 222.210 51.560 ;
        RECT 222.455 51.480 222.760 51.940 ;
        RECT 222.930 51.230 223.185 51.760 ;
        RECT 223.420 51.480 223.665 51.940 ;
        RECT 221.890 51.030 222.215 51.205 ;
        RECT 221.890 50.730 222.805 51.030 ;
        RECT 222.065 50.700 222.805 50.730 ;
        RECT 219.540 50.370 220.215 50.530 ;
        RECT 220.675 50.450 220.845 50.540 ;
        RECT 219.540 50.360 220.505 50.370 ;
        RECT 219.180 50.190 219.350 50.330 ;
        RECT 215.925 49.390 216.175 49.850 ;
        RECT 216.345 49.560 216.595 49.890 ;
        RECT 216.810 49.560 217.490 49.890 ;
        RECT 217.660 49.990 218.735 50.160 ;
        RECT 219.180 50.020 219.740 50.190 ;
        RECT 220.045 50.070 220.505 50.360 ;
        RECT 220.675 50.280 221.895 50.450 ;
        RECT 217.660 49.650 217.830 49.990 ;
        RECT 218.065 49.390 218.395 49.820 ;
        RECT 218.565 49.650 218.735 49.990 ;
        RECT 219.030 49.390 219.400 49.850 ;
        RECT 219.570 49.560 219.740 50.020 ;
        RECT 220.675 49.900 220.845 50.280 ;
        RECT 222.065 50.110 222.235 50.700 ;
        RECT 222.975 50.580 223.185 51.230 ;
        RECT 223.360 50.700 223.675 51.310 ;
        RECT 223.845 50.950 224.095 51.760 ;
        RECT 224.265 51.415 224.525 51.940 ;
        RECT 224.695 51.290 224.955 51.745 ;
        RECT 225.125 51.460 225.385 51.940 ;
        RECT 225.555 51.290 225.815 51.745 ;
        RECT 225.985 51.460 226.245 51.940 ;
        RECT 226.415 51.290 226.675 51.745 ;
        RECT 226.845 51.460 227.105 51.940 ;
        RECT 227.275 51.290 227.535 51.745 ;
        RECT 227.705 51.460 228.005 51.940 ;
        RECT 224.695 51.120 228.005 51.290 ;
        RECT 223.845 50.700 226.865 50.950 ;
        RECT 219.975 49.560 220.845 49.900 ;
        RECT 221.435 49.940 222.235 50.110 ;
        RECT 221.015 49.390 221.265 49.850 ;
        RECT 221.435 49.650 221.605 49.940 ;
        RECT 221.785 49.390 222.115 49.770 ;
        RECT 222.455 49.390 222.760 50.530 ;
        RECT 222.930 49.700 223.185 50.580 ;
        RECT 223.370 49.390 223.665 50.500 ;
        RECT 223.845 49.565 224.095 50.700 ;
        RECT 227.035 50.530 228.005 51.120 ;
        RECT 228.420 51.170 230.090 51.940 ;
        RECT 230.265 51.390 230.520 51.680 ;
        RECT 230.690 51.560 231.020 51.940 ;
        RECT 230.265 51.220 231.015 51.390 ;
        RECT 228.420 50.650 229.170 51.170 ;
        RECT 224.265 49.390 224.525 50.500 ;
        RECT 224.695 50.290 228.005 50.530 ;
        RECT 229.340 50.480 230.090 51.000 ;
        RECT 224.695 49.565 224.955 50.290 ;
        RECT 225.125 49.390 225.385 50.120 ;
        RECT 225.555 49.565 225.815 50.290 ;
        RECT 225.985 49.390 226.245 50.120 ;
        RECT 226.415 49.565 226.675 50.290 ;
        RECT 226.845 49.390 227.105 50.120 ;
        RECT 227.275 49.565 227.535 50.290 ;
        RECT 227.705 49.390 228.000 50.120 ;
        RECT 228.420 49.390 230.090 50.480 ;
        RECT 230.265 50.400 230.615 51.050 ;
        RECT 230.785 50.230 231.015 51.220 ;
        RECT 230.265 50.060 231.015 50.230 ;
        RECT 230.265 49.560 230.520 50.060 ;
        RECT 230.690 49.390 231.020 49.890 ;
        RECT 231.190 49.560 231.360 51.680 ;
        RECT 231.720 51.580 232.050 51.940 ;
        RECT 232.220 51.550 232.715 51.720 ;
        RECT 232.920 51.550 233.775 51.720 ;
        RECT 231.590 50.360 232.050 51.410 ;
        RECT 231.530 49.575 231.855 50.360 ;
        RECT 232.220 50.190 232.390 51.550 ;
        RECT 232.560 50.640 232.910 51.260 ;
        RECT 233.080 51.040 233.435 51.260 ;
        RECT 233.080 50.450 233.250 51.040 ;
        RECT 233.605 50.840 233.775 51.550 ;
        RECT 234.650 51.480 234.980 51.940 ;
        RECT 235.190 51.580 235.540 51.750 ;
        RECT 233.980 51.010 234.770 51.260 ;
        RECT 235.190 51.190 235.450 51.580 ;
        RECT 235.760 51.490 236.710 51.770 ;
        RECT 236.880 51.500 237.070 51.940 ;
        RECT 237.240 51.560 238.310 51.730 ;
        RECT 234.940 50.840 235.110 51.020 ;
        RECT 232.220 50.020 232.615 50.190 ;
        RECT 232.785 50.060 233.250 50.450 ;
        RECT 233.420 50.670 235.110 50.840 ;
        RECT 232.445 49.890 232.615 50.020 ;
        RECT 233.420 49.890 233.590 50.670 ;
        RECT 235.280 50.500 235.450 51.190 ;
        RECT 233.950 50.330 235.450 50.500 ;
        RECT 235.640 50.530 235.850 51.320 ;
        RECT 236.020 50.700 236.370 51.320 ;
        RECT 236.540 50.710 236.710 51.490 ;
        RECT 237.240 51.330 237.410 51.560 ;
        RECT 236.880 51.160 237.410 51.330 ;
        RECT 236.880 50.880 237.100 51.160 ;
        RECT 237.580 50.990 237.820 51.390 ;
        RECT 236.540 50.540 236.945 50.710 ;
        RECT 237.280 50.620 237.820 50.990 ;
        RECT 237.990 51.205 238.310 51.560 ;
        RECT 238.555 51.480 238.860 51.940 ;
        RECT 239.030 51.230 239.285 51.760 ;
        RECT 237.990 51.030 238.315 51.205 ;
        RECT 237.990 50.730 238.905 51.030 ;
        RECT 238.165 50.700 238.905 50.730 ;
        RECT 235.640 50.370 236.315 50.530 ;
        RECT 236.775 50.450 236.945 50.540 ;
        RECT 235.640 50.360 236.605 50.370 ;
        RECT 235.280 50.190 235.450 50.330 ;
        RECT 232.025 49.390 232.275 49.850 ;
        RECT 232.445 49.560 232.695 49.890 ;
        RECT 232.910 49.560 233.590 49.890 ;
        RECT 233.760 49.990 234.835 50.160 ;
        RECT 235.280 50.020 235.840 50.190 ;
        RECT 236.145 50.070 236.605 50.360 ;
        RECT 236.775 50.280 237.995 50.450 ;
        RECT 233.760 49.650 233.930 49.990 ;
        RECT 234.165 49.390 234.495 49.820 ;
        RECT 234.665 49.650 234.835 49.990 ;
        RECT 235.130 49.390 235.500 49.850 ;
        RECT 235.670 49.560 235.840 50.020 ;
        RECT 236.775 49.900 236.945 50.280 ;
        RECT 238.165 50.110 238.335 50.700 ;
        RECT 239.075 50.580 239.285 51.230 ;
        RECT 239.460 51.215 239.750 51.940 ;
        RECT 236.075 49.560 236.945 49.900 ;
        RECT 237.535 49.940 238.335 50.110 ;
        RECT 237.115 49.390 237.365 49.850 ;
        RECT 237.535 49.650 237.705 49.940 ;
        RECT 237.885 49.390 238.215 49.770 ;
        RECT 238.555 49.390 238.860 50.530 ;
        RECT 239.030 49.700 239.285 50.580 ;
        RECT 239.920 51.120 240.605 51.760 ;
        RECT 240.775 51.120 240.945 51.940 ;
        RECT 241.115 51.290 241.445 51.755 ;
        RECT 241.615 51.470 241.785 51.940 ;
        RECT 242.045 51.550 243.230 51.720 ;
        RECT 243.400 51.380 243.730 51.770 ;
        RECT 242.430 51.290 242.815 51.380 ;
        RECT 241.115 51.120 242.815 51.290 ;
        RECT 243.220 51.200 243.730 51.380 ;
        RECT 239.460 49.390 239.750 50.555 ;
        RECT 239.920 50.150 240.170 51.120 ;
        RECT 240.340 50.740 240.675 50.950 ;
        RECT 240.845 50.740 241.295 50.950 ;
        RECT 241.485 50.920 241.970 50.950 ;
        RECT 241.485 50.750 241.990 50.920 ;
        RECT 241.485 50.740 241.970 50.750 ;
        RECT 240.505 50.570 240.675 50.740 ;
        RECT 240.505 50.400 241.425 50.570 ;
        RECT 239.920 49.560 240.585 50.150 ;
        RECT 240.755 49.390 241.085 50.230 ;
        RECT 241.255 50.150 241.425 50.400 ;
        RECT 241.595 50.320 241.970 50.740 ;
        RECT 242.160 50.700 242.540 50.950 ;
        RECT 242.720 50.740 243.050 50.950 ;
        RECT 242.160 50.320 242.480 50.700 ;
        RECT 243.220 50.570 243.390 51.200 ;
        RECT 244.060 51.170 246.650 51.940 ;
        RECT 243.560 50.740 243.890 51.030 ;
        RECT 244.060 50.650 245.270 51.170 ;
        RECT 246.820 51.120 247.505 51.760 ;
        RECT 247.675 51.120 247.845 51.940 ;
        RECT 248.015 51.290 248.345 51.755 ;
        RECT 248.515 51.470 248.685 51.940 ;
        RECT 248.945 51.550 250.130 51.720 ;
        RECT 250.300 51.380 250.630 51.770 ;
        RECT 249.330 51.290 249.715 51.380 ;
        RECT 248.015 51.120 249.715 51.290 ;
        RECT 250.120 51.200 250.630 51.380 ;
        RECT 250.960 51.200 251.345 51.770 ;
        RECT 251.515 51.480 251.840 51.940 ;
        RECT 252.360 51.310 252.640 51.770 ;
        RECT 242.650 50.400 243.735 50.570 ;
        RECT 245.440 50.480 246.650 51.000 ;
        RECT 242.650 50.150 242.820 50.400 ;
        RECT 241.255 49.980 242.820 50.150 ;
        RECT 241.595 49.560 242.400 49.980 ;
        RECT 242.990 49.390 243.240 50.230 ;
        RECT 243.435 49.560 243.735 50.400 ;
        RECT 244.060 49.390 246.650 50.480 ;
        RECT 246.820 50.150 247.070 51.120 ;
        RECT 247.240 50.740 247.575 50.950 ;
        RECT 247.745 50.740 248.195 50.950 ;
        RECT 248.385 50.920 248.870 50.950 ;
        RECT 248.385 50.750 248.890 50.920 ;
        RECT 248.385 50.740 248.870 50.750 ;
        RECT 247.405 50.570 247.575 50.740 ;
        RECT 247.405 50.400 248.325 50.570 ;
        RECT 246.820 49.560 247.485 50.150 ;
        RECT 247.655 49.390 247.985 50.230 ;
        RECT 248.155 50.150 248.325 50.400 ;
        RECT 248.495 50.320 248.870 50.740 ;
        RECT 249.060 50.700 249.440 50.950 ;
        RECT 249.620 50.740 249.950 50.950 ;
        RECT 249.060 50.320 249.380 50.700 ;
        RECT 250.120 50.570 250.290 51.200 ;
        RECT 250.460 50.740 250.790 51.030 ;
        RECT 249.550 50.400 250.635 50.570 ;
        RECT 249.550 50.150 249.720 50.400 ;
        RECT 248.155 49.980 249.720 50.150 ;
        RECT 248.495 49.560 249.300 49.980 ;
        RECT 249.890 49.390 250.140 50.230 ;
        RECT 250.335 49.560 250.635 50.400 ;
        RECT 250.960 50.530 251.240 51.200 ;
        RECT 251.515 51.140 252.640 51.310 ;
        RECT 251.515 51.030 251.965 51.140 ;
        RECT 251.410 50.700 251.965 51.030 ;
        RECT 252.830 50.970 253.230 51.770 ;
        RECT 253.630 51.480 253.900 51.940 ;
        RECT 254.070 51.310 254.355 51.770 ;
        RECT 250.960 49.560 251.345 50.530 ;
        RECT 251.515 50.240 251.965 50.700 ;
        RECT 252.135 50.410 253.230 50.970 ;
        RECT 251.515 50.020 252.640 50.240 ;
        RECT 251.515 49.390 251.840 49.850 ;
        RECT 252.360 49.560 252.640 50.020 ;
        RECT 252.830 49.560 253.230 50.410 ;
        RECT 253.400 51.140 254.355 51.310 ;
        RECT 254.640 51.190 255.850 51.940 ;
        RECT 256.025 51.390 256.280 51.680 ;
        RECT 256.450 51.560 256.780 51.940 ;
        RECT 256.025 51.220 256.775 51.390 ;
        RECT 253.400 50.240 253.610 51.140 ;
        RECT 253.780 50.410 254.470 50.970 ;
        RECT 254.640 50.650 255.160 51.190 ;
        RECT 255.330 50.480 255.850 51.020 ;
        RECT 253.400 50.020 254.355 50.240 ;
        RECT 253.630 49.390 253.900 49.850 ;
        RECT 254.070 49.560 254.355 50.020 ;
        RECT 254.640 49.390 255.850 50.480 ;
        RECT 256.025 50.400 256.375 51.050 ;
        RECT 256.545 50.230 256.775 51.220 ;
        RECT 256.025 50.060 256.775 50.230 ;
        RECT 256.025 49.560 256.280 50.060 ;
        RECT 256.450 49.390 256.780 49.890 ;
        RECT 256.950 49.560 257.120 51.680 ;
        RECT 257.480 51.580 257.810 51.940 ;
        RECT 257.980 51.550 258.475 51.720 ;
        RECT 258.680 51.550 259.535 51.720 ;
        RECT 257.350 50.360 257.810 51.410 ;
        RECT 257.290 49.575 257.615 50.360 ;
        RECT 257.980 50.190 258.150 51.550 ;
        RECT 258.320 50.640 258.670 51.260 ;
        RECT 258.840 51.040 259.195 51.260 ;
        RECT 258.840 50.450 259.010 51.040 ;
        RECT 259.365 50.840 259.535 51.550 ;
        RECT 260.410 51.480 260.740 51.940 ;
        RECT 260.950 51.580 261.300 51.750 ;
        RECT 259.740 51.010 260.530 51.260 ;
        RECT 260.950 51.190 261.210 51.580 ;
        RECT 261.520 51.490 262.470 51.770 ;
        RECT 262.640 51.500 262.830 51.940 ;
        RECT 263.000 51.560 264.070 51.730 ;
        RECT 260.700 50.840 260.870 51.020 ;
        RECT 257.980 50.020 258.375 50.190 ;
        RECT 258.545 50.060 259.010 50.450 ;
        RECT 259.180 50.670 260.870 50.840 ;
        RECT 258.205 49.890 258.375 50.020 ;
        RECT 259.180 49.890 259.350 50.670 ;
        RECT 261.040 50.500 261.210 51.190 ;
        RECT 259.710 50.330 261.210 50.500 ;
        RECT 261.400 50.530 261.610 51.320 ;
        RECT 261.780 50.700 262.130 51.320 ;
        RECT 262.300 50.710 262.470 51.490 ;
        RECT 263.000 51.330 263.170 51.560 ;
        RECT 262.640 51.160 263.170 51.330 ;
        RECT 262.640 50.880 262.860 51.160 ;
        RECT 263.340 50.990 263.580 51.390 ;
        RECT 262.300 50.540 262.705 50.710 ;
        RECT 263.040 50.620 263.580 50.990 ;
        RECT 263.750 51.205 264.070 51.560 ;
        RECT 264.315 51.480 264.620 51.940 ;
        RECT 264.790 51.230 265.045 51.760 ;
        RECT 263.750 51.030 264.075 51.205 ;
        RECT 263.750 50.730 264.665 51.030 ;
        RECT 263.925 50.700 264.665 50.730 ;
        RECT 261.400 50.370 262.075 50.530 ;
        RECT 262.535 50.450 262.705 50.540 ;
        RECT 261.400 50.360 262.365 50.370 ;
        RECT 261.040 50.190 261.210 50.330 ;
        RECT 257.785 49.390 258.035 49.850 ;
        RECT 258.205 49.560 258.455 49.890 ;
        RECT 258.670 49.560 259.350 49.890 ;
        RECT 259.520 49.990 260.595 50.160 ;
        RECT 261.040 50.020 261.600 50.190 ;
        RECT 261.905 50.070 262.365 50.360 ;
        RECT 262.535 50.280 263.755 50.450 ;
        RECT 259.520 49.650 259.690 49.990 ;
        RECT 259.925 49.390 260.255 49.820 ;
        RECT 260.425 49.650 260.595 49.990 ;
        RECT 260.890 49.390 261.260 49.850 ;
        RECT 261.430 49.560 261.600 50.020 ;
        RECT 262.535 49.900 262.705 50.280 ;
        RECT 263.925 50.110 264.095 50.700 ;
        RECT 264.835 50.580 265.045 51.230 ;
        RECT 265.220 51.215 265.510 51.940 ;
        RECT 265.680 51.170 267.350 51.940 ;
        RECT 267.985 51.390 268.240 51.680 ;
        RECT 268.410 51.560 268.740 51.940 ;
        RECT 267.985 51.220 268.735 51.390 ;
        RECT 265.680 50.650 266.430 51.170 ;
        RECT 261.835 49.560 262.705 49.900 ;
        RECT 263.295 49.940 264.095 50.110 ;
        RECT 262.875 49.390 263.125 49.850 ;
        RECT 263.295 49.650 263.465 49.940 ;
        RECT 263.645 49.390 263.975 49.770 ;
        RECT 264.315 49.390 264.620 50.530 ;
        RECT 264.790 49.700 265.045 50.580 ;
        RECT 265.220 49.390 265.510 50.555 ;
        RECT 266.600 50.480 267.350 51.000 ;
        RECT 265.680 49.390 267.350 50.480 ;
        RECT 267.985 50.400 268.335 51.050 ;
        RECT 268.505 50.230 268.735 51.220 ;
        RECT 267.985 50.060 268.735 50.230 ;
        RECT 267.985 49.560 268.240 50.060 ;
        RECT 268.410 49.390 268.740 49.890 ;
        RECT 268.910 49.560 269.080 51.680 ;
        RECT 269.440 51.580 269.770 51.940 ;
        RECT 269.940 51.550 270.435 51.720 ;
        RECT 270.640 51.550 271.495 51.720 ;
        RECT 269.310 50.360 269.770 51.410 ;
        RECT 269.250 49.575 269.575 50.360 ;
        RECT 269.940 50.190 270.110 51.550 ;
        RECT 270.280 50.640 270.630 51.260 ;
        RECT 270.800 51.040 271.155 51.260 ;
        RECT 270.800 50.450 270.970 51.040 ;
        RECT 271.325 50.840 271.495 51.550 ;
        RECT 272.370 51.480 272.700 51.940 ;
        RECT 272.910 51.580 273.260 51.750 ;
        RECT 271.700 51.010 272.490 51.260 ;
        RECT 272.910 51.190 273.170 51.580 ;
        RECT 273.480 51.490 274.430 51.770 ;
        RECT 274.600 51.500 274.790 51.940 ;
        RECT 274.960 51.560 276.030 51.730 ;
        RECT 272.660 50.840 272.830 51.020 ;
        RECT 269.940 50.020 270.335 50.190 ;
        RECT 270.505 50.060 270.970 50.450 ;
        RECT 271.140 50.670 272.830 50.840 ;
        RECT 270.165 49.890 270.335 50.020 ;
        RECT 271.140 49.890 271.310 50.670 ;
        RECT 273.000 50.500 273.170 51.190 ;
        RECT 271.670 50.330 273.170 50.500 ;
        RECT 273.360 50.530 273.570 51.320 ;
        RECT 273.740 50.700 274.090 51.320 ;
        RECT 274.260 50.710 274.430 51.490 ;
        RECT 274.960 51.330 275.130 51.560 ;
        RECT 274.600 51.160 275.130 51.330 ;
        RECT 274.600 50.880 274.820 51.160 ;
        RECT 275.300 50.990 275.540 51.390 ;
        RECT 274.260 50.540 274.665 50.710 ;
        RECT 275.000 50.620 275.540 50.990 ;
        RECT 275.710 51.205 276.030 51.560 ;
        RECT 276.275 51.480 276.580 51.940 ;
        RECT 276.750 51.230 277.005 51.760 ;
        RECT 275.710 51.030 276.035 51.205 ;
        RECT 275.710 50.730 276.625 51.030 ;
        RECT 275.885 50.700 276.625 50.730 ;
        RECT 273.360 50.370 274.035 50.530 ;
        RECT 274.495 50.450 274.665 50.540 ;
        RECT 273.360 50.360 274.325 50.370 ;
        RECT 273.000 50.190 273.170 50.330 ;
        RECT 269.745 49.390 269.995 49.850 ;
        RECT 270.165 49.560 270.415 49.890 ;
        RECT 270.630 49.560 271.310 49.890 ;
        RECT 271.480 49.990 272.555 50.160 ;
        RECT 273.000 50.020 273.560 50.190 ;
        RECT 273.865 50.070 274.325 50.360 ;
        RECT 274.495 50.280 275.715 50.450 ;
        RECT 271.480 49.650 271.650 49.990 ;
        RECT 271.885 49.390 272.215 49.820 ;
        RECT 272.385 49.650 272.555 49.990 ;
        RECT 272.850 49.390 273.220 49.850 ;
        RECT 273.390 49.560 273.560 50.020 ;
        RECT 274.495 49.900 274.665 50.280 ;
        RECT 275.885 50.110 276.055 50.700 ;
        RECT 276.795 50.580 277.005 51.230 ;
        RECT 273.795 49.560 274.665 49.900 ;
        RECT 275.255 49.940 276.055 50.110 ;
        RECT 274.835 49.390 275.085 49.850 ;
        RECT 275.255 49.650 275.425 49.940 ;
        RECT 275.605 49.390 275.935 49.770 ;
        RECT 276.275 49.390 276.580 50.530 ;
        RECT 276.750 49.700 277.005 50.580 ;
        RECT 277.185 51.230 277.440 51.760 ;
        RECT 277.610 51.480 277.915 51.940 ;
        RECT 278.160 51.560 279.230 51.730 ;
        RECT 277.185 50.580 277.395 51.230 ;
        RECT 278.160 51.205 278.480 51.560 ;
        RECT 278.155 51.030 278.480 51.205 ;
        RECT 277.565 50.730 278.480 51.030 ;
        RECT 278.650 50.990 278.890 51.390 ;
        RECT 279.060 51.330 279.230 51.560 ;
        RECT 279.400 51.500 279.590 51.940 ;
        RECT 279.760 51.490 280.710 51.770 ;
        RECT 280.930 51.580 281.280 51.750 ;
        RECT 279.060 51.160 279.590 51.330 ;
        RECT 277.565 50.700 278.305 50.730 ;
        RECT 277.185 49.700 277.440 50.580 ;
        RECT 277.610 49.390 277.915 50.530 ;
        RECT 278.135 50.110 278.305 50.700 ;
        RECT 278.650 50.620 279.190 50.990 ;
        RECT 279.370 50.880 279.590 51.160 ;
        RECT 279.760 50.710 279.930 51.490 ;
        RECT 279.525 50.540 279.930 50.710 ;
        RECT 280.100 50.700 280.450 51.320 ;
        RECT 279.525 50.450 279.695 50.540 ;
        RECT 280.620 50.530 280.830 51.320 ;
        RECT 278.475 50.280 279.695 50.450 ;
        RECT 280.155 50.370 280.830 50.530 ;
        RECT 278.135 49.940 278.935 50.110 ;
        RECT 278.255 49.390 278.585 49.770 ;
        RECT 278.765 49.650 278.935 49.940 ;
        RECT 279.525 49.900 279.695 50.280 ;
        RECT 279.865 50.360 280.830 50.370 ;
        RECT 281.020 51.190 281.280 51.580 ;
        RECT 281.490 51.480 281.820 51.940 ;
        RECT 282.695 51.550 283.550 51.720 ;
        RECT 283.755 51.550 284.250 51.720 ;
        RECT 284.420 51.580 284.750 51.940 ;
        RECT 281.020 50.500 281.190 51.190 ;
        RECT 281.360 50.840 281.530 51.020 ;
        RECT 281.700 51.010 282.490 51.260 ;
        RECT 282.695 50.840 282.865 51.550 ;
        RECT 283.035 51.040 283.390 51.260 ;
        RECT 281.360 50.670 283.050 50.840 ;
        RECT 279.865 50.070 280.325 50.360 ;
        RECT 281.020 50.330 282.520 50.500 ;
        RECT 281.020 50.190 281.190 50.330 ;
        RECT 280.630 50.020 281.190 50.190 ;
        RECT 279.105 49.390 279.355 49.850 ;
        RECT 279.525 49.560 280.395 49.900 ;
        RECT 280.630 49.560 280.800 50.020 ;
        RECT 281.635 49.990 282.710 50.160 ;
        RECT 280.970 49.390 281.340 49.850 ;
        RECT 281.635 49.650 281.805 49.990 ;
        RECT 281.975 49.390 282.305 49.820 ;
        RECT 282.540 49.650 282.710 49.990 ;
        RECT 282.880 49.890 283.050 50.670 ;
        RECT 283.220 50.450 283.390 51.040 ;
        RECT 283.560 50.640 283.910 51.260 ;
        RECT 283.220 50.060 283.685 50.450 ;
        RECT 284.080 50.190 284.250 51.550 ;
        RECT 284.420 50.360 284.880 51.410 ;
        RECT 283.855 50.020 284.250 50.190 ;
        RECT 283.855 49.890 284.025 50.020 ;
        RECT 282.880 49.560 283.560 49.890 ;
        RECT 283.775 49.560 284.025 49.890 ;
        RECT 284.195 49.390 284.445 49.850 ;
        RECT 284.615 49.575 284.940 50.360 ;
        RECT 285.110 49.560 285.280 51.680 ;
        RECT 285.450 51.560 285.780 51.940 ;
        RECT 285.950 51.390 286.205 51.680 ;
        RECT 285.455 51.220 286.205 51.390 ;
        RECT 285.455 50.230 285.685 51.220 ;
        RECT 286.380 51.200 286.765 51.770 ;
        RECT 286.935 51.480 287.260 51.940 ;
        RECT 287.780 51.310 288.060 51.770 ;
        RECT 285.855 50.400 286.205 51.050 ;
        RECT 286.380 50.530 286.660 51.200 ;
        RECT 286.935 51.140 288.060 51.310 ;
        RECT 286.935 51.030 287.385 51.140 ;
        RECT 286.830 50.700 287.385 51.030 ;
        RECT 288.250 50.970 288.650 51.770 ;
        RECT 289.050 51.480 289.320 51.940 ;
        RECT 289.490 51.310 289.775 51.770 ;
        RECT 285.455 50.060 286.205 50.230 ;
        RECT 285.450 49.390 285.780 49.890 ;
        RECT 285.950 49.560 286.205 50.060 ;
        RECT 286.380 49.560 286.765 50.530 ;
        RECT 286.935 50.240 287.385 50.700 ;
        RECT 287.555 50.410 288.650 50.970 ;
        RECT 286.935 50.020 288.060 50.240 ;
        RECT 286.935 49.390 287.260 49.850 ;
        RECT 287.780 49.560 288.060 50.020 ;
        RECT 288.250 49.560 288.650 50.410 ;
        RECT 288.820 51.140 289.775 51.310 ;
        RECT 290.980 51.215 291.270 51.940 ;
        RECT 291.920 51.470 292.215 51.940 ;
        RECT 292.385 51.300 292.645 51.745 ;
        RECT 292.815 51.470 293.075 51.940 ;
        RECT 293.245 51.300 293.500 51.745 ;
        RECT 293.670 51.470 293.970 51.940 ;
        RECT 288.820 50.240 289.030 51.140 ;
        RECT 291.460 51.130 294.490 51.300 ;
        RECT 289.200 50.410 289.890 50.970 ;
        RECT 291.460 50.565 291.630 51.130 ;
        RECT 291.800 50.735 294.015 50.960 ;
        RECT 294.190 50.565 294.490 51.130 ;
        RECT 294.660 51.170 298.170 51.940 ;
        RECT 298.340 51.190 299.550 51.940 ;
        RECT 300.095 51.600 300.350 51.760 ;
        RECT 300.010 51.430 300.350 51.600 ;
        RECT 300.530 51.480 300.815 51.940 ;
        RECT 300.095 51.230 300.350 51.430 ;
        RECT 294.660 50.650 296.310 51.170 ;
        RECT 288.820 50.020 289.775 50.240 ;
        RECT 289.050 49.390 289.320 49.850 ;
        RECT 289.490 49.560 289.775 50.020 ;
        RECT 290.980 49.390 291.270 50.555 ;
        RECT 291.460 50.395 294.490 50.565 ;
        RECT 296.480 50.480 298.170 51.000 ;
        RECT 298.340 50.650 298.860 51.190 ;
        RECT 299.030 50.480 299.550 51.020 ;
        RECT 291.440 49.390 291.785 50.225 ;
        RECT 291.960 49.590 292.215 50.395 ;
        RECT 292.385 49.390 292.645 50.225 ;
        RECT 292.820 49.590 293.075 50.395 ;
        RECT 293.245 49.390 293.505 50.225 ;
        RECT 293.675 49.590 293.935 50.395 ;
        RECT 294.105 49.390 294.490 50.225 ;
        RECT 294.660 49.390 298.170 50.480 ;
        RECT 298.340 49.390 299.550 50.480 ;
        RECT 300.095 50.370 300.275 51.230 ;
        RECT 300.995 51.030 301.245 51.680 ;
        RECT 300.445 50.700 301.245 51.030 ;
        RECT 300.095 49.700 300.350 50.370 ;
        RECT 300.530 49.390 300.815 50.190 ;
        RECT 300.995 50.110 301.245 50.700 ;
        RECT 301.445 51.345 301.765 51.675 ;
        RECT 301.945 51.460 302.605 51.940 ;
        RECT 302.805 51.550 303.655 51.720 ;
        RECT 301.445 50.450 301.635 51.345 ;
        RECT 301.955 51.020 302.615 51.290 ;
        RECT 302.285 50.960 302.615 51.020 ;
        RECT 301.805 50.790 302.135 50.850 ;
        RECT 302.805 50.790 302.975 51.550 ;
        RECT 304.215 51.480 304.535 51.940 ;
        RECT 304.735 51.300 304.985 51.730 ;
        RECT 305.275 51.500 305.685 51.940 ;
        RECT 305.855 51.560 306.870 51.760 ;
        RECT 303.145 51.130 304.395 51.300 ;
        RECT 303.145 51.010 303.475 51.130 ;
        RECT 301.805 50.620 303.705 50.790 ;
        RECT 301.445 50.280 303.365 50.450 ;
        RECT 301.445 50.260 301.765 50.280 ;
        RECT 300.995 49.600 301.325 50.110 ;
        RECT 301.595 49.650 301.765 50.260 ;
        RECT 303.535 50.110 303.705 50.620 ;
        RECT 303.875 50.550 304.055 50.960 ;
        RECT 304.225 50.370 304.395 51.130 ;
        RECT 301.935 49.390 302.265 50.080 ;
        RECT 302.495 49.940 303.705 50.110 ;
        RECT 303.875 50.060 304.395 50.370 ;
        RECT 304.565 50.960 304.985 51.300 ;
        RECT 305.275 50.960 305.685 51.290 ;
        RECT 304.565 50.190 304.755 50.960 ;
        RECT 305.855 50.830 306.025 51.560 ;
        RECT 307.170 51.390 307.340 51.720 ;
        RECT 307.510 51.560 307.840 51.940 ;
        RECT 306.195 51.010 306.545 51.380 ;
        RECT 305.855 50.790 306.275 50.830 ;
        RECT 304.925 50.620 306.275 50.790 ;
        RECT 304.925 50.460 305.175 50.620 ;
        RECT 305.685 50.190 305.935 50.450 ;
        RECT 304.565 49.940 305.935 50.190 ;
        RECT 302.495 49.650 302.735 49.940 ;
        RECT 303.535 49.860 303.705 49.940 ;
        RECT 302.935 49.390 303.355 49.770 ;
        RECT 303.535 49.610 304.165 49.860 ;
        RECT 304.635 49.390 304.965 49.770 ;
        RECT 305.135 49.650 305.305 49.940 ;
        RECT 306.105 49.775 306.275 50.620 ;
        RECT 306.725 50.450 306.945 51.320 ;
        RECT 307.170 51.200 307.865 51.390 ;
        RECT 306.445 50.070 306.945 50.450 ;
        RECT 307.115 50.400 307.525 51.020 ;
        RECT 307.695 50.230 307.865 51.200 ;
        RECT 307.170 50.060 307.865 50.230 ;
        RECT 305.485 49.390 305.865 49.770 ;
        RECT 306.105 49.605 306.935 49.775 ;
        RECT 307.170 49.560 307.340 50.060 ;
        RECT 307.510 49.390 307.840 49.890 ;
        RECT 308.055 49.560 308.280 51.680 ;
        RECT 308.450 51.560 308.780 51.940 ;
        RECT 308.950 51.390 309.120 51.680 ;
        RECT 308.455 51.220 309.120 51.390 ;
        RECT 308.455 50.230 308.685 51.220 ;
        RECT 309.840 51.190 311.050 51.940 ;
        RECT 308.855 50.400 309.205 51.050 ;
        RECT 309.840 50.480 310.360 51.020 ;
        RECT 310.530 50.650 311.050 51.190 ;
        RECT 308.455 50.060 309.120 50.230 ;
        RECT 308.450 49.390 308.780 49.890 ;
        RECT 308.950 49.560 309.120 50.060 ;
        RECT 309.840 49.390 311.050 50.480 ;
        RECT 162.095 49.220 311.135 49.390 ;
        RECT 162.180 48.130 163.390 49.220 ;
        RECT 163.560 48.785 168.905 49.220 ;
        RECT 169.080 48.785 174.425 49.220 ;
        RECT 162.180 47.420 162.700 47.960 ;
        RECT 162.870 47.590 163.390 48.130 ;
        RECT 162.180 46.670 163.390 47.420 ;
        RECT 165.145 47.215 165.485 48.045 ;
        RECT 166.965 47.535 167.315 48.785 ;
        RECT 170.665 47.215 171.005 48.045 ;
        RECT 172.485 47.535 172.835 48.785 ;
        RECT 175.060 48.055 175.350 49.220 ;
        RECT 175.525 48.080 175.860 49.050 ;
        RECT 176.030 48.080 176.200 49.220 ;
        RECT 176.370 48.880 178.400 49.050 ;
        RECT 175.525 47.410 175.695 48.080 ;
        RECT 176.370 47.910 176.540 48.880 ;
        RECT 175.865 47.580 176.120 47.910 ;
        RECT 176.345 47.580 176.540 47.910 ;
        RECT 176.710 48.540 177.835 48.710 ;
        RECT 175.950 47.410 176.120 47.580 ;
        RECT 176.710 47.410 176.880 48.540 ;
        RECT 163.560 46.670 168.905 47.215 ;
        RECT 169.080 46.670 174.425 47.215 ;
        RECT 175.060 46.670 175.350 47.395 ;
        RECT 175.525 46.840 175.780 47.410 ;
        RECT 175.950 47.240 176.880 47.410 ;
        RECT 177.050 48.200 178.060 48.370 ;
        RECT 177.050 47.400 177.220 48.200 ;
        RECT 177.425 47.520 177.700 48.000 ;
        RECT 177.420 47.350 177.700 47.520 ;
        RECT 176.705 47.205 176.880 47.240 ;
        RECT 175.950 46.670 176.280 47.070 ;
        RECT 176.705 46.840 177.235 47.205 ;
        RECT 177.425 46.840 177.700 47.350 ;
        RECT 177.870 46.840 178.060 48.200 ;
        RECT 178.230 48.215 178.400 48.880 ;
        RECT 178.570 48.460 178.740 49.220 ;
        RECT 178.975 48.460 179.490 48.870 ;
        RECT 178.230 48.025 178.980 48.215 ;
        RECT 179.150 47.650 179.490 48.460 ;
        RECT 178.260 47.480 179.490 47.650 ;
        RECT 179.665 48.080 180.000 49.050 ;
        RECT 180.170 48.080 180.340 49.220 ;
        RECT 180.510 48.880 182.540 49.050 ;
        RECT 178.240 46.670 178.750 47.205 ;
        RECT 178.970 46.875 179.215 47.480 ;
        RECT 179.665 47.410 179.835 48.080 ;
        RECT 180.510 47.910 180.680 48.880 ;
        RECT 180.005 47.580 180.260 47.910 ;
        RECT 180.485 47.580 180.680 47.910 ;
        RECT 180.850 48.540 181.975 48.710 ;
        RECT 180.090 47.410 180.260 47.580 ;
        RECT 180.850 47.410 181.020 48.540 ;
        RECT 179.665 46.840 179.920 47.410 ;
        RECT 180.090 47.240 181.020 47.410 ;
        RECT 181.190 48.200 182.200 48.370 ;
        RECT 181.190 47.400 181.360 48.200 ;
        RECT 180.845 47.205 181.020 47.240 ;
        RECT 180.090 46.670 180.420 47.070 ;
        RECT 180.845 46.840 181.375 47.205 ;
        RECT 181.565 47.180 181.840 48.000 ;
        RECT 181.560 47.010 181.840 47.180 ;
        RECT 181.565 46.840 181.840 47.010 ;
        RECT 182.010 46.840 182.200 48.200 ;
        RECT 182.370 48.215 182.540 48.880 ;
        RECT 182.710 48.460 182.880 49.220 ;
        RECT 183.115 48.460 183.630 48.870 ;
        RECT 182.370 48.025 183.120 48.215 ;
        RECT 183.290 47.650 183.630 48.460 ;
        RECT 184.270 48.080 184.600 49.220 ;
        RECT 185.130 48.250 185.460 49.035 ;
        RECT 184.780 48.080 185.460 48.250 ;
        RECT 185.640 48.130 188.230 49.220 ;
        RECT 184.260 47.660 184.610 47.910 ;
        RECT 182.400 47.480 183.630 47.650 ;
        RECT 184.780 47.480 184.950 48.080 ;
        RECT 185.120 47.660 185.470 47.910 ;
        RECT 182.380 46.670 182.890 47.205 ;
        RECT 183.110 46.875 183.355 47.480 ;
        RECT 184.270 46.670 184.540 47.480 ;
        RECT 184.710 46.840 185.040 47.480 ;
        RECT 185.210 46.670 185.450 47.480 ;
        RECT 185.640 47.440 186.850 47.960 ;
        RECT 187.020 47.610 188.230 48.130 ;
        RECT 188.440 48.080 188.670 49.220 ;
        RECT 188.840 48.070 189.170 49.050 ;
        RECT 189.340 48.080 189.550 49.220 ;
        RECT 189.780 48.130 193.290 49.220 ;
        RECT 193.460 48.130 194.670 49.220 ;
        RECT 195.090 48.490 195.385 49.220 ;
        RECT 195.555 48.320 195.815 49.045 ;
        RECT 195.985 48.490 196.245 49.220 ;
        RECT 196.415 48.320 196.675 49.045 ;
        RECT 196.845 48.490 197.105 49.220 ;
        RECT 197.275 48.320 197.535 49.045 ;
        RECT 197.705 48.490 197.965 49.220 ;
        RECT 198.135 48.320 198.395 49.045 ;
        RECT 188.420 47.660 188.750 47.910 ;
        RECT 185.640 46.670 188.230 47.440 ;
        RECT 188.440 46.670 188.670 47.490 ;
        RECT 188.920 47.470 189.170 48.070 ;
        RECT 188.840 46.840 189.170 47.470 ;
        RECT 189.340 46.670 189.550 47.490 ;
        RECT 189.780 47.440 191.430 47.960 ;
        RECT 191.600 47.610 193.290 48.130 ;
        RECT 189.780 46.670 193.290 47.440 ;
        RECT 193.460 47.420 193.980 47.960 ;
        RECT 194.150 47.590 194.670 48.130 ;
        RECT 195.085 48.080 198.395 48.320 ;
        RECT 198.565 48.110 198.825 49.220 ;
        RECT 195.085 47.490 196.055 48.080 ;
        RECT 198.995 47.910 199.245 49.045 ;
        RECT 199.425 48.110 199.720 49.220 ;
        RECT 200.820 48.055 201.110 49.220 ;
        RECT 201.280 48.785 206.625 49.220 ;
        RECT 206.800 48.785 212.145 49.220 ;
        RECT 196.225 47.660 199.245 47.910 ;
        RECT 193.460 46.670 194.670 47.420 ;
        RECT 195.085 47.320 198.395 47.490 ;
        RECT 195.085 46.670 195.385 47.150 ;
        RECT 195.555 46.865 195.815 47.320 ;
        RECT 195.985 46.670 196.245 47.150 ;
        RECT 196.415 46.865 196.675 47.320 ;
        RECT 196.845 46.670 197.105 47.150 ;
        RECT 197.275 46.865 197.535 47.320 ;
        RECT 197.705 46.670 197.965 47.150 ;
        RECT 198.135 46.865 198.395 47.320 ;
        RECT 198.565 46.670 198.825 47.195 ;
        RECT 198.995 46.850 199.245 47.660 ;
        RECT 199.415 47.300 199.730 47.910 ;
        RECT 199.425 46.670 199.670 47.130 ;
        RECT 200.820 46.670 201.110 47.395 ;
        RECT 202.865 47.215 203.205 48.045 ;
        RECT 204.685 47.535 205.035 48.785 ;
        RECT 208.385 47.215 208.725 48.045 ;
        RECT 210.205 47.535 210.555 48.785 ;
        RECT 212.320 48.130 213.990 49.220 ;
        RECT 212.320 47.440 213.070 47.960 ;
        RECT 213.240 47.610 213.990 48.130 ;
        RECT 214.195 48.430 214.730 49.050 ;
        RECT 201.280 46.670 206.625 47.215 ;
        RECT 206.800 46.670 212.145 47.215 ;
        RECT 212.320 46.670 213.990 47.440 ;
        RECT 214.195 47.410 214.510 48.430 ;
        RECT 214.900 48.420 215.230 49.220 ;
        RECT 216.465 48.550 216.720 49.050 ;
        RECT 216.890 48.720 217.220 49.220 ;
        RECT 215.715 48.250 216.105 48.425 ;
        RECT 216.465 48.380 217.215 48.550 ;
        RECT 214.680 48.080 216.105 48.250 ;
        RECT 214.680 47.580 214.850 48.080 ;
        RECT 214.195 46.840 214.810 47.410 ;
        RECT 215.100 47.350 215.365 47.910 ;
        RECT 215.535 47.180 215.705 48.080 ;
        RECT 215.875 47.350 216.230 47.910 ;
        RECT 216.465 47.560 216.815 48.210 ;
        RECT 216.985 47.390 217.215 48.380 ;
        RECT 216.465 47.220 217.215 47.390 ;
        RECT 214.980 46.670 215.195 47.180 ;
        RECT 215.425 46.850 215.705 47.180 ;
        RECT 215.885 46.670 216.125 47.180 ;
        RECT 216.465 46.930 216.720 47.220 ;
        RECT 216.890 46.670 217.220 47.050 ;
        RECT 217.390 46.930 217.560 49.050 ;
        RECT 217.730 48.250 218.055 49.035 ;
        RECT 218.225 48.760 218.475 49.220 ;
        RECT 218.645 48.720 218.895 49.050 ;
        RECT 219.110 48.720 219.790 49.050 ;
        RECT 218.645 48.590 218.815 48.720 ;
        RECT 218.420 48.420 218.815 48.590 ;
        RECT 217.790 47.200 218.250 48.250 ;
        RECT 218.420 47.060 218.590 48.420 ;
        RECT 218.985 48.160 219.450 48.550 ;
        RECT 218.760 47.350 219.110 47.970 ;
        RECT 219.280 47.570 219.450 48.160 ;
        RECT 219.620 47.940 219.790 48.720 ;
        RECT 219.960 48.620 220.130 48.960 ;
        RECT 220.365 48.790 220.695 49.220 ;
        RECT 220.865 48.620 221.035 48.960 ;
        RECT 221.330 48.760 221.700 49.220 ;
        RECT 219.960 48.450 221.035 48.620 ;
        RECT 221.870 48.590 222.040 49.050 ;
        RECT 222.275 48.710 223.145 49.050 ;
        RECT 223.315 48.760 223.565 49.220 ;
        RECT 221.480 48.420 222.040 48.590 ;
        RECT 221.480 48.280 221.650 48.420 ;
        RECT 220.150 48.110 221.650 48.280 ;
        RECT 222.345 48.250 222.805 48.540 ;
        RECT 219.620 47.770 221.310 47.940 ;
        RECT 219.280 47.350 219.635 47.570 ;
        RECT 219.805 47.060 219.975 47.770 ;
        RECT 220.180 47.350 220.970 47.600 ;
        RECT 221.140 47.590 221.310 47.770 ;
        RECT 221.480 47.420 221.650 48.110 ;
        RECT 217.920 46.670 218.250 47.030 ;
        RECT 218.420 46.890 218.915 47.060 ;
        RECT 219.120 46.890 219.975 47.060 ;
        RECT 220.850 46.670 221.180 47.130 ;
        RECT 221.390 47.030 221.650 47.420 ;
        RECT 221.840 48.240 222.805 48.250 ;
        RECT 222.975 48.330 223.145 48.710 ;
        RECT 223.735 48.670 223.905 48.960 ;
        RECT 224.085 48.840 224.415 49.220 ;
        RECT 223.735 48.500 224.535 48.670 ;
        RECT 221.840 48.080 222.515 48.240 ;
        RECT 222.975 48.160 224.195 48.330 ;
        RECT 221.840 47.290 222.050 48.080 ;
        RECT 222.975 48.070 223.145 48.160 ;
        RECT 222.220 47.290 222.570 47.910 ;
        RECT 222.740 47.900 223.145 48.070 ;
        RECT 222.740 47.120 222.910 47.900 ;
        RECT 223.080 47.450 223.300 47.730 ;
        RECT 223.480 47.620 224.020 47.990 ;
        RECT 224.365 47.910 224.535 48.500 ;
        RECT 224.755 48.080 225.060 49.220 ;
        RECT 225.230 48.030 225.485 48.910 ;
        RECT 226.580 48.055 226.870 49.220 ;
        RECT 227.040 48.130 228.250 49.220 ;
        RECT 228.535 48.590 228.820 49.050 ;
        RECT 228.990 48.760 229.260 49.220 ;
        RECT 228.535 48.370 229.490 48.590 ;
        RECT 224.365 47.880 225.105 47.910 ;
        RECT 223.080 47.280 223.610 47.450 ;
        RECT 221.390 46.860 221.740 47.030 ;
        RECT 221.960 46.840 222.910 47.120 ;
        RECT 223.080 46.670 223.270 47.110 ;
        RECT 223.440 47.050 223.610 47.280 ;
        RECT 223.780 47.220 224.020 47.620 ;
        RECT 224.190 47.580 225.105 47.880 ;
        RECT 224.190 47.405 224.515 47.580 ;
        RECT 224.190 47.050 224.510 47.405 ;
        RECT 225.275 47.380 225.485 48.030 ;
        RECT 227.040 47.420 227.560 47.960 ;
        RECT 227.730 47.590 228.250 48.130 ;
        RECT 228.420 47.640 229.110 48.200 ;
        RECT 229.280 47.470 229.490 48.370 ;
        RECT 223.440 46.880 224.510 47.050 ;
        RECT 224.755 46.670 225.060 47.130 ;
        RECT 225.230 46.850 225.485 47.380 ;
        RECT 226.580 46.670 226.870 47.395 ;
        RECT 227.040 46.670 228.250 47.420 ;
        RECT 228.535 47.300 229.490 47.470 ;
        RECT 229.660 48.200 230.060 49.050 ;
        RECT 230.250 48.590 230.530 49.050 ;
        RECT 231.050 48.760 231.375 49.220 ;
        RECT 230.250 48.370 231.375 48.590 ;
        RECT 229.660 47.640 230.755 48.200 ;
        RECT 230.925 47.910 231.375 48.370 ;
        RECT 231.545 48.080 231.930 49.050 ;
        RECT 232.105 48.550 232.360 49.050 ;
        RECT 232.530 48.720 232.860 49.220 ;
        RECT 232.105 48.380 232.855 48.550 ;
        RECT 228.535 46.840 228.820 47.300 ;
        RECT 228.990 46.670 229.260 47.130 ;
        RECT 229.660 46.840 230.060 47.640 ;
        RECT 230.925 47.580 231.480 47.910 ;
        RECT 230.925 47.470 231.375 47.580 ;
        RECT 230.250 47.300 231.375 47.470 ;
        RECT 231.650 47.410 231.930 48.080 ;
        RECT 232.105 47.560 232.455 48.210 ;
        RECT 230.250 46.840 230.530 47.300 ;
        RECT 231.050 46.670 231.375 47.130 ;
        RECT 231.545 46.840 231.930 47.410 ;
        RECT 232.625 47.390 232.855 48.380 ;
        RECT 232.105 47.220 232.855 47.390 ;
        RECT 232.105 46.930 232.360 47.220 ;
        RECT 232.530 46.670 232.860 47.050 ;
        RECT 233.030 46.930 233.200 49.050 ;
        RECT 233.370 48.250 233.695 49.035 ;
        RECT 233.865 48.760 234.115 49.220 ;
        RECT 234.285 48.720 234.535 49.050 ;
        RECT 234.750 48.720 235.430 49.050 ;
        RECT 234.285 48.590 234.455 48.720 ;
        RECT 234.060 48.420 234.455 48.590 ;
        RECT 233.430 47.200 233.890 48.250 ;
        RECT 234.060 47.060 234.230 48.420 ;
        RECT 234.625 48.160 235.090 48.550 ;
        RECT 234.400 47.350 234.750 47.970 ;
        RECT 234.920 47.570 235.090 48.160 ;
        RECT 235.260 47.940 235.430 48.720 ;
        RECT 235.600 48.620 235.770 48.960 ;
        RECT 236.005 48.790 236.335 49.220 ;
        RECT 236.505 48.620 236.675 48.960 ;
        RECT 236.970 48.760 237.340 49.220 ;
        RECT 235.600 48.450 236.675 48.620 ;
        RECT 237.510 48.590 237.680 49.050 ;
        RECT 237.915 48.710 238.785 49.050 ;
        RECT 238.955 48.760 239.205 49.220 ;
        RECT 237.120 48.420 237.680 48.590 ;
        RECT 237.120 48.280 237.290 48.420 ;
        RECT 235.790 48.110 237.290 48.280 ;
        RECT 237.985 48.250 238.445 48.540 ;
        RECT 235.260 47.770 236.950 47.940 ;
        RECT 234.920 47.350 235.275 47.570 ;
        RECT 235.445 47.060 235.615 47.770 ;
        RECT 235.820 47.350 236.610 47.600 ;
        RECT 236.780 47.590 236.950 47.770 ;
        RECT 237.120 47.420 237.290 48.110 ;
        RECT 233.560 46.670 233.890 47.030 ;
        RECT 234.060 46.890 234.555 47.060 ;
        RECT 234.760 46.890 235.615 47.060 ;
        RECT 236.490 46.670 236.820 47.130 ;
        RECT 237.030 47.030 237.290 47.420 ;
        RECT 237.480 48.240 238.445 48.250 ;
        RECT 238.615 48.330 238.785 48.710 ;
        RECT 239.375 48.670 239.545 48.960 ;
        RECT 239.725 48.840 240.055 49.220 ;
        RECT 239.375 48.500 240.175 48.670 ;
        RECT 237.480 48.080 238.155 48.240 ;
        RECT 238.615 48.160 239.835 48.330 ;
        RECT 237.480 47.290 237.690 48.080 ;
        RECT 238.615 48.070 238.785 48.160 ;
        RECT 237.860 47.290 238.210 47.910 ;
        RECT 238.380 47.900 238.785 48.070 ;
        RECT 238.380 47.120 238.550 47.900 ;
        RECT 238.720 47.450 238.940 47.730 ;
        RECT 239.120 47.620 239.660 47.990 ;
        RECT 240.005 47.910 240.175 48.500 ;
        RECT 240.395 48.080 240.700 49.220 ;
        RECT 240.870 48.030 241.125 48.910 ;
        RECT 240.005 47.880 240.745 47.910 ;
        RECT 238.720 47.280 239.250 47.450 ;
        RECT 237.030 46.860 237.380 47.030 ;
        RECT 237.600 46.840 238.550 47.120 ;
        RECT 238.720 46.670 238.910 47.110 ;
        RECT 239.080 47.050 239.250 47.280 ;
        RECT 239.420 47.220 239.660 47.620 ;
        RECT 239.830 47.580 240.745 47.880 ;
        RECT 239.830 47.405 240.155 47.580 ;
        RECT 239.830 47.050 240.150 47.405 ;
        RECT 240.915 47.380 241.125 48.030 ;
        RECT 239.080 46.880 240.150 47.050 ;
        RECT 240.395 46.670 240.700 47.130 ;
        RECT 240.870 46.850 241.125 47.380 ;
        RECT 241.305 48.030 241.560 48.910 ;
        RECT 241.730 48.080 242.035 49.220 ;
        RECT 242.375 48.840 242.705 49.220 ;
        RECT 242.885 48.670 243.055 48.960 ;
        RECT 243.225 48.760 243.475 49.220 ;
        RECT 242.255 48.500 243.055 48.670 ;
        RECT 243.645 48.710 244.515 49.050 ;
        RECT 241.305 47.380 241.515 48.030 ;
        RECT 242.255 47.910 242.425 48.500 ;
        RECT 243.645 48.330 243.815 48.710 ;
        RECT 244.750 48.590 244.920 49.050 ;
        RECT 245.090 48.760 245.460 49.220 ;
        RECT 245.755 48.620 245.925 48.960 ;
        RECT 246.095 48.790 246.425 49.220 ;
        RECT 246.660 48.620 246.830 48.960 ;
        RECT 242.595 48.160 243.815 48.330 ;
        RECT 243.985 48.250 244.445 48.540 ;
        RECT 244.750 48.420 245.310 48.590 ;
        RECT 245.755 48.450 246.830 48.620 ;
        RECT 247.000 48.720 247.680 49.050 ;
        RECT 247.895 48.720 248.145 49.050 ;
        RECT 248.315 48.760 248.565 49.220 ;
        RECT 245.140 48.280 245.310 48.420 ;
        RECT 243.985 48.240 244.950 48.250 ;
        RECT 243.645 48.070 243.815 48.160 ;
        RECT 244.275 48.080 244.950 48.240 ;
        RECT 241.685 47.880 242.425 47.910 ;
        RECT 241.685 47.580 242.600 47.880 ;
        RECT 242.275 47.405 242.600 47.580 ;
        RECT 241.305 46.850 241.560 47.380 ;
        RECT 241.730 46.670 242.035 47.130 ;
        RECT 242.280 47.050 242.600 47.405 ;
        RECT 242.770 47.620 243.310 47.990 ;
        RECT 243.645 47.900 244.050 48.070 ;
        RECT 242.770 47.220 243.010 47.620 ;
        RECT 243.490 47.450 243.710 47.730 ;
        RECT 243.180 47.280 243.710 47.450 ;
        RECT 243.180 47.050 243.350 47.280 ;
        RECT 243.880 47.120 244.050 47.900 ;
        RECT 244.220 47.290 244.570 47.910 ;
        RECT 244.740 47.290 244.950 48.080 ;
        RECT 245.140 48.110 246.640 48.280 ;
        RECT 245.140 47.420 245.310 48.110 ;
        RECT 247.000 47.940 247.170 48.720 ;
        RECT 247.975 48.590 248.145 48.720 ;
        RECT 245.480 47.770 247.170 47.940 ;
        RECT 247.340 48.160 247.805 48.550 ;
        RECT 247.975 48.420 248.370 48.590 ;
        RECT 245.480 47.590 245.650 47.770 ;
        RECT 242.280 46.880 243.350 47.050 ;
        RECT 243.520 46.670 243.710 47.110 ;
        RECT 243.880 46.840 244.830 47.120 ;
        RECT 245.140 47.030 245.400 47.420 ;
        RECT 245.820 47.350 246.610 47.600 ;
        RECT 245.050 46.860 245.400 47.030 ;
        RECT 245.610 46.670 245.940 47.130 ;
        RECT 246.815 47.060 246.985 47.770 ;
        RECT 247.340 47.570 247.510 48.160 ;
        RECT 247.155 47.350 247.510 47.570 ;
        RECT 247.680 47.350 248.030 47.970 ;
        RECT 248.200 47.060 248.370 48.420 ;
        RECT 248.735 48.250 249.060 49.035 ;
        RECT 248.540 47.200 249.000 48.250 ;
        RECT 246.815 46.890 247.670 47.060 ;
        RECT 247.875 46.890 248.370 47.060 ;
        RECT 248.540 46.670 248.870 47.030 ;
        RECT 249.230 46.930 249.400 49.050 ;
        RECT 249.570 48.720 249.900 49.220 ;
        RECT 250.070 48.550 250.325 49.050 ;
        RECT 249.575 48.380 250.325 48.550 ;
        RECT 249.575 47.390 249.805 48.380 ;
        RECT 249.975 47.560 250.325 48.210 ;
        RECT 250.500 48.130 252.170 49.220 ;
        RECT 250.500 47.440 251.250 47.960 ;
        RECT 251.420 47.610 252.170 48.130 ;
        RECT 252.340 48.055 252.630 49.220 ;
        RECT 252.845 48.080 253.140 49.220 ;
        RECT 253.400 48.250 253.730 49.050 ;
        RECT 253.900 48.420 254.070 49.220 ;
        RECT 254.240 48.250 254.570 49.050 ;
        RECT 254.740 48.420 254.910 49.220 ;
        RECT 255.080 48.270 255.410 49.050 ;
        RECT 255.580 48.760 255.750 49.220 ;
        RECT 256.025 48.550 256.280 49.050 ;
        RECT 256.450 48.720 256.780 49.220 ;
        RECT 256.025 48.380 256.775 48.550 ;
        RECT 255.080 48.250 255.850 48.270 ;
        RECT 253.400 48.080 255.850 48.250 ;
        RECT 252.820 47.660 255.330 47.910 ;
        RECT 255.500 47.490 255.850 48.080 ;
        RECT 256.025 47.560 256.375 48.210 ;
        RECT 249.575 47.220 250.325 47.390 ;
        RECT 249.570 46.670 249.900 47.050 ;
        RECT 250.070 46.930 250.325 47.220 ;
        RECT 250.500 46.670 252.170 47.440 ;
        RECT 252.340 46.670 252.630 47.395 ;
        RECT 253.480 47.310 255.850 47.490 ;
        RECT 256.545 47.390 256.775 48.380 ;
        RECT 252.845 46.670 253.110 47.130 ;
        RECT 253.480 46.840 253.650 47.310 ;
        RECT 253.900 46.670 254.070 47.130 ;
        RECT 254.320 46.840 254.490 47.310 ;
        RECT 254.740 46.670 254.910 47.130 ;
        RECT 255.160 46.840 255.330 47.310 ;
        RECT 256.025 47.220 256.775 47.390 ;
        RECT 255.500 46.670 255.750 47.135 ;
        RECT 256.025 46.930 256.280 47.220 ;
        RECT 256.450 46.670 256.780 47.050 ;
        RECT 256.950 46.930 257.120 49.050 ;
        RECT 257.290 48.250 257.615 49.035 ;
        RECT 257.785 48.760 258.035 49.220 ;
        RECT 258.205 48.720 258.455 49.050 ;
        RECT 258.670 48.720 259.350 49.050 ;
        RECT 258.205 48.590 258.375 48.720 ;
        RECT 257.980 48.420 258.375 48.590 ;
        RECT 257.350 47.200 257.810 48.250 ;
        RECT 257.980 47.060 258.150 48.420 ;
        RECT 258.545 48.160 259.010 48.550 ;
        RECT 258.320 47.350 258.670 47.970 ;
        RECT 258.840 47.570 259.010 48.160 ;
        RECT 259.180 47.940 259.350 48.720 ;
        RECT 259.520 48.620 259.690 48.960 ;
        RECT 259.925 48.790 260.255 49.220 ;
        RECT 260.425 48.620 260.595 48.960 ;
        RECT 260.890 48.760 261.260 49.220 ;
        RECT 259.520 48.450 260.595 48.620 ;
        RECT 261.430 48.590 261.600 49.050 ;
        RECT 261.835 48.710 262.705 49.050 ;
        RECT 262.875 48.760 263.125 49.220 ;
        RECT 261.040 48.420 261.600 48.590 ;
        RECT 261.040 48.280 261.210 48.420 ;
        RECT 259.710 48.110 261.210 48.280 ;
        RECT 261.905 48.250 262.365 48.540 ;
        RECT 259.180 47.770 260.870 47.940 ;
        RECT 258.840 47.350 259.195 47.570 ;
        RECT 259.365 47.060 259.535 47.770 ;
        RECT 259.740 47.350 260.530 47.600 ;
        RECT 260.700 47.590 260.870 47.770 ;
        RECT 261.040 47.420 261.210 48.110 ;
        RECT 257.480 46.670 257.810 47.030 ;
        RECT 257.980 46.890 258.475 47.060 ;
        RECT 258.680 46.890 259.535 47.060 ;
        RECT 260.410 46.670 260.740 47.130 ;
        RECT 260.950 47.030 261.210 47.420 ;
        RECT 261.400 48.240 262.365 48.250 ;
        RECT 262.535 48.330 262.705 48.710 ;
        RECT 263.295 48.670 263.465 48.960 ;
        RECT 263.645 48.840 263.975 49.220 ;
        RECT 263.295 48.500 264.095 48.670 ;
        RECT 261.400 48.080 262.075 48.240 ;
        RECT 262.535 48.160 263.755 48.330 ;
        RECT 261.400 47.290 261.610 48.080 ;
        RECT 262.535 48.070 262.705 48.160 ;
        RECT 261.780 47.290 262.130 47.910 ;
        RECT 262.300 47.900 262.705 48.070 ;
        RECT 262.300 47.120 262.470 47.900 ;
        RECT 262.640 47.450 262.860 47.730 ;
        RECT 263.040 47.620 263.580 47.990 ;
        RECT 263.925 47.910 264.095 48.500 ;
        RECT 264.315 48.080 264.620 49.220 ;
        RECT 264.790 48.030 265.045 48.910 ;
        RECT 265.220 48.665 265.825 49.220 ;
        RECT 266.000 48.710 266.480 49.050 ;
        RECT 266.650 48.675 266.905 49.220 ;
        RECT 265.220 48.565 265.835 48.665 ;
        RECT 265.650 48.540 265.835 48.565 ;
        RECT 263.925 47.880 264.665 47.910 ;
        RECT 262.640 47.280 263.170 47.450 ;
        RECT 260.950 46.860 261.300 47.030 ;
        RECT 261.520 46.840 262.470 47.120 ;
        RECT 262.640 46.670 262.830 47.110 ;
        RECT 263.000 47.050 263.170 47.280 ;
        RECT 263.340 47.220 263.580 47.620 ;
        RECT 263.750 47.580 264.665 47.880 ;
        RECT 263.750 47.405 264.075 47.580 ;
        RECT 263.750 47.050 264.070 47.405 ;
        RECT 264.835 47.380 265.045 48.030 ;
        RECT 265.220 47.945 265.480 48.395 ;
        RECT 265.650 48.295 265.980 48.540 ;
        RECT 266.150 48.220 266.905 48.470 ;
        RECT 267.075 48.350 267.350 49.050 ;
        RECT 267.625 48.760 267.795 49.220 ;
        RECT 267.965 48.590 268.295 49.050 ;
        RECT 266.135 48.185 266.905 48.220 ;
        RECT 266.120 48.175 266.905 48.185 ;
        RECT 266.115 48.160 267.010 48.175 ;
        RECT 266.095 48.145 267.010 48.160 ;
        RECT 266.075 48.135 267.010 48.145 ;
        RECT 266.050 48.125 267.010 48.135 ;
        RECT 265.980 48.095 267.010 48.125 ;
        RECT 265.960 48.065 267.010 48.095 ;
        RECT 265.940 48.035 267.010 48.065 ;
        RECT 265.910 48.010 267.010 48.035 ;
        RECT 265.875 47.975 267.010 48.010 ;
        RECT 265.845 47.970 267.010 47.975 ;
        RECT 265.845 47.965 266.235 47.970 ;
        RECT 265.845 47.955 266.210 47.965 ;
        RECT 265.845 47.950 266.195 47.955 ;
        RECT 265.845 47.945 266.180 47.950 ;
        RECT 265.220 47.940 266.180 47.945 ;
        RECT 265.220 47.930 266.170 47.940 ;
        RECT 265.220 47.925 266.160 47.930 ;
        RECT 265.220 47.915 266.150 47.925 ;
        RECT 265.220 47.905 266.145 47.915 ;
        RECT 265.220 47.900 266.140 47.905 ;
        RECT 265.220 47.885 266.130 47.900 ;
        RECT 265.220 47.870 266.125 47.885 ;
        RECT 265.220 47.845 266.115 47.870 ;
        RECT 265.220 47.775 266.110 47.845 ;
        RECT 263.000 46.880 264.070 47.050 ;
        RECT 264.315 46.670 264.620 47.130 ;
        RECT 264.790 46.850 265.045 47.380 ;
        RECT 265.220 47.220 265.770 47.605 ;
        RECT 265.940 47.050 266.110 47.775 ;
        RECT 265.220 46.880 266.110 47.050 ;
        RECT 266.280 47.375 266.610 47.800 ;
        RECT 266.780 47.575 267.010 47.970 ;
        RECT 266.280 47.350 266.530 47.375 ;
        RECT 266.280 46.890 266.500 47.350 ;
        RECT 267.180 47.320 267.350 48.350 ;
        RECT 266.670 46.670 266.920 47.210 ;
        RECT 267.090 46.840 267.350 47.320 ;
        RECT 267.520 48.420 268.295 48.590 ;
        RECT 268.465 48.420 268.635 49.220 ;
        RECT 267.520 47.410 267.950 48.420 ;
        RECT 269.220 48.250 269.580 48.425 ;
        RECT 269.925 48.420 270.180 49.220 ;
        RECT 270.350 48.250 270.680 49.050 ;
        RECT 270.850 48.420 271.020 49.220 ;
        RECT 271.190 48.250 271.520 49.050 ;
        RECT 268.120 48.080 269.580 48.250 ;
        RECT 269.820 48.080 271.520 48.250 ;
        RECT 271.690 48.080 271.950 49.220 ;
        RECT 272.120 48.785 277.465 49.220 ;
        RECT 268.120 47.580 268.290 48.080 ;
        RECT 267.520 47.240 268.215 47.410 ;
        RECT 268.460 47.350 268.870 47.910 ;
        RECT 267.545 46.670 267.875 47.070 ;
        RECT 268.045 46.970 268.215 47.240 ;
        RECT 269.040 47.180 269.220 48.080 ;
        RECT 269.390 47.860 269.585 47.910 ;
        RECT 269.390 47.690 269.590 47.860 ;
        RECT 269.390 47.350 269.585 47.690 ;
        RECT 269.820 47.490 270.100 48.080 ;
        RECT 270.270 47.660 271.020 47.910 ;
        RECT 271.190 47.660 271.950 47.910 ;
        RECT 269.820 47.240 270.680 47.490 ;
        RECT 270.850 47.300 271.950 47.470 ;
        RECT 268.385 46.670 268.700 47.180 ;
        RECT 268.930 46.840 269.220 47.180 ;
        RECT 269.390 46.670 269.630 47.180 ;
        RECT 269.930 47.050 270.260 47.070 ;
        RECT 270.850 47.050 271.100 47.300 ;
        RECT 269.930 46.840 271.100 47.050 ;
        RECT 271.270 46.670 271.440 47.130 ;
        RECT 271.610 46.840 271.950 47.300 ;
        RECT 273.705 47.215 274.045 48.045 ;
        RECT 275.525 47.535 275.875 48.785 ;
        RECT 278.100 48.055 278.390 49.220 ;
        RECT 278.560 48.460 279.075 48.870 ;
        RECT 279.310 48.460 279.480 49.220 ;
        RECT 279.650 48.880 281.680 49.050 ;
        RECT 278.560 47.650 278.900 48.460 ;
        RECT 279.650 48.215 279.820 48.880 ;
        RECT 280.215 48.540 281.340 48.710 ;
        RECT 279.070 48.025 279.820 48.215 ;
        RECT 279.990 48.200 281.000 48.370 ;
        RECT 278.560 47.480 279.790 47.650 ;
        RECT 272.120 46.670 277.465 47.215 ;
        RECT 278.100 46.670 278.390 47.395 ;
        RECT 278.835 46.875 279.080 47.480 ;
        RECT 279.300 46.670 279.810 47.205 ;
        RECT 279.990 46.840 280.180 48.200 ;
        RECT 280.350 47.860 280.625 48.000 ;
        RECT 280.350 47.690 280.630 47.860 ;
        RECT 280.350 46.840 280.625 47.690 ;
        RECT 280.830 47.400 281.000 48.200 ;
        RECT 281.170 47.410 281.340 48.540 ;
        RECT 281.510 47.910 281.680 48.880 ;
        RECT 281.850 48.080 282.020 49.220 ;
        RECT 282.190 48.080 282.525 49.050 ;
        RECT 283.625 48.550 283.880 49.050 ;
        RECT 284.050 48.720 284.380 49.220 ;
        RECT 283.625 48.380 284.375 48.550 ;
        RECT 281.510 47.580 281.705 47.910 ;
        RECT 281.930 47.580 282.185 47.910 ;
        RECT 281.930 47.410 282.100 47.580 ;
        RECT 282.355 47.410 282.525 48.080 ;
        RECT 283.625 47.560 283.975 48.210 ;
        RECT 281.170 47.240 282.100 47.410 ;
        RECT 281.170 47.205 281.345 47.240 ;
        RECT 280.815 46.840 281.345 47.205 ;
        RECT 281.770 46.670 282.100 47.070 ;
        RECT 282.270 46.840 282.525 47.410 ;
        RECT 284.145 47.390 284.375 48.380 ;
        RECT 283.625 47.220 284.375 47.390 ;
        RECT 283.625 46.930 283.880 47.220 ;
        RECT 284.050 46.670 284.380 47.050 ;
        RECT 284.550 46.930 284.720 49.050 ;
        RECT 284.890 48.250 285.215 49.035 ;
        RECT 285.385 48.760 285.635 49.220 ;
        RECT 285.805 48.720 286.055 49.050 ;
        RECT 286.270 48.720 286.950 49.050 ;
        RECT 285.805 48.590 285.975 48.720 ;
        RECT 285.580 48.420 285.975 48.590 ;
        RECT 284.950 47.200 285.410 48.250 ;
        RECT 285.580 47.060 285.750 48.420 ;
        RECT 286.145 48.160 286.610 48.550 ;
        RECT 285.920 47.350 286.270 47.970 ;
        RECT 286.440 47.570 286.610 48.160 ;
        RECT 286.780 47.940 286.950 48.720 ;
        RECT 287.120 48.620 287.290 48.960 ;
        RECT 287.525 48.790 287.855 49.220 ;
        RECT 288.025 48.620 288.195 48.960 ;
        RECT 288.490 48.760 288.860 49.220 ;
        RECT 287.120 48.450 288.195 48.620 ;
        RECT 289.030 48.590 289.200 49.050 ;
        RECT 289.435 48.710 290.305 49.050 ;
        RECT 290.475 48.760 290.725 49.220 ;
        RECT 288.640 48.420 289.200 48.590 ;
        RECT 288.640 48.280 288.810 48.420 ;
        RECT 287.310 48.110 288.810 48.280 ;
        RECT 289.505 48.250 289.965 48.540 ;
        RECT 286.780 47.770 288.470 47.940 ;
        RECT 286.440 47.350 286.795 47.570 ;
        RECT 286.965 47.060 287.135 47.770 ;
        RECT 287.340 47.350 288.130 47.600 ;
        RECT 288.300 47.590 288.470 47.770 ;
        RECT 288.640 47.420 288.810 48.110 ;
        RECT 285.080 46.670 285.410 47.030 ;
        RECT 285.580 46.890 286.075 47.060 ;
        RECT 286.280 46.890 287.135 47.060 ;
        RECT 288.010 46.670 288.340 47.130 ;
        RECT 288.550 47.030 288.810 47.420 ;
        RECT 289.000 48.240 289.965 48.250 ;
        RECT 290.135 48.330 290.305 48.710 ;
        RECT 290.895 48.670 291.065 48.960 ;
        RECT 291.245 48.840 291.575 49.220 ;
        RECT 290.895 48.500 291.695 48.670 ;
        RECT 289.000 48.080 289.675 48.240 ;
        RECT 290.135 48.160 291.355 48.330 ;
        RECT 289.000 47.290 289.210 48.080 ;
        RECT 290.135 48.070 290.305 48.160 ;
        RECT 289.380 47.290 289.730 47.910 ;
        RECT 289.900 47.900 290.305 48.070 ;
        RECT 289.900 47.120 290.070 47.900 ;
        RECT 290.240 47.450 290.460 47.730 ;
        RECT 290.640 47.620 291.180 47.990 ;
        RECT 291.525 47.910 291.695 48.500 ;
        RECT 291.915 48.080 292.220 49.220 ;
        RECT 292.390 48.030 292.645 48.910 ;
        RECT 291.525 47.880 292.265 47.910 ;
        RECT 290.240 47.280 290.770 47.450 ;
        RECT 288.550 46.860 288.900 47.030 ;
        RECT 289.120 46.840 290.070 47.120 ;
        RECT 290.240 46.670 290.430 47.110 ;
        RECT 290.600 47.050 290.770 47.280 ;
        RECT 290.940 47.220 291.180 47.620 ;
        RECT 291.350 47.580 292.265 47.880 ;
        RECT 291.350 47.405 291.675 47.580 ;
        RECT 291.350 47.050 291.670 47.405 ;
        RECT 292.435 47.380 292.645 48.030 ;
        RECT 290.600 46.880 291.670 47.050 ;
        RECT 291.915 46.670 292.220 47.130 ;
        RECT 292.390 46.850 292.645 47.380 ;
        RECT 292.820 48.080 293.205 49.050 ;
        RECT 293.375 48.760 293.700 49.220 ;
        RECT 294.220 48.590 294.500 49.050 ;
        RECT 293.375 48.370 294.500 48.590 ;
        RECT 292.820 47.410 293.100 48.080 ;
        RECT 293.375 47.910 293.825 48.370 ;
        RECT 294.690 48.200 295.090 49.050 ;
        RECT 295.490 48.760 295.760 49.220 ;
        RECT 295.930 48.590 296.215 49.050 ;
        RECT 296.500 48.785 301.845 49.220 ;
        RECT 293.270 47.580 293.825 47.910 ;
        RECT 293.995 47.640 295.090 48.200 ;
        RECT 293.375 47.470 293.825 47.580 ;
        RECT 292.820 46.840 293.205 47.410 ;
        RECT 293.375 47.300 294.500 47.470 ;
        RECT 293.375 46.670 293.700 47.130 ;
        RECT 294.220 46.840 294.500 47.300 ;
        RECT 294.690 46.840 295.090 47.640 ;
        RECT 295.260 48.370 296.215 48.590 ;
        RECT 295.260 47.470 295.470 48.370 ;
        RECT 295.640 47.640 296.330 48.200 ;
        RECT 295.260 47.300 296.215 47.470 ;
        RECT 295.490 46.670 295.760 47.130 ;
        RECT 295.930 46.840 296.215 47.300 ;
        RECT 298.085 47.215 298.425 48.045 ;
        RECT 299.905 47.535 300.255 48.785 ;
        RECT 302.020 48.130 303.690 49.220 ;
        RECT 302.020 47.440 302.770 47.960 ;
        RECT 302.940 47.610 303.690 48.130 ;
        RECT 303.860 48.055 304.150 49.220 ;
        RECT 304.320 48.785 309.665 49.220 ;
        RECT 296.500 46.670 301.845 47.215 ;
        RECT 302.020 46.670 303.690 47.440 ;
        RECT 303.860 46.670 304.150 47.395 ;
        RECT 305.905 47.215 306.245 48.045 ;
        RECT 307.725 47.535 308.075 48.785 ;
        RECT 309.840 48.130 311.050 49.220 ;
        RECT 309.840 47.590 310.360 48.130 ;
        RECT 310.530 47.420 311.050 47.960 ;
        RECT 304.320 46.670 309.665 47.215 ;
        RECT 309.840 46.670 311.050 47.420 ;
        RECT 162.095 46.500 311.135 46.670 ;
        RECT 162.180 45.750 163.390 46.500 ;
        RECT 163.560 45.955 168.905 46.500 ;
        RECT 162.180 45.210 162.700 45.750 ;
        RECT 162.870 45.040 163.390 45.580 ;
        RECT 165.145 45.125 165.485 45.955 ;
        RECT 169.080 45.730 172.590 46.500 ;
        RECT 172.765 45.950 173.020 46.240 ;
        RECT 173.190 46.120 173.520 46.500 ;
        RECT 172.765 45.780 173.515 45.950 ;
        RECT 162.180 43.950 163.390 45.040 ;
        RECT 166.965 44.385 167.315 45.635 ;
        RECT 169.080 45.210 170.730 45.730 ;
        RECT 170.900 45.040 172.590 45.560 ;
        RECT 163.560 43.950 168.905 44.385 ;
        RECT 169.080 43.950 172.590 45.040 ;
        RECT 172.765 44.960 173.115 45.610 ;
        RECT 173.285 44.790 173.515 45.780 ;
        RECT 172.765 44.620 173.515 44.790 ;
        RECT 172.765 44.120 173.020 44.620 ;
        RECT 173.190 43.950 173.520 44.450 ;
        RECT 173.690 44.120 173.860 46.240 ;
        RECT 174.220 46.140 174.550 46.500 ;
        RECT 174.720 46.110 175.215 46.280 ;
        RECT 175.420 46.110 176.275 46.280 ;
        RECT 174.090 44.920 174.550 45.970 ;
        RECT 174.030 44.135 174.355 44.920 ;
        RECT 174.720 44.750 174.890 46.110 ;
        RECT 175.060 45.200 175.410 45.820 ;
        RECT 175.580 45.600 175.935 45.820 ;
        RECT 175.580 45.010 175.750 45.600 ;
        RECT 176.105 45.400 176.275 46.110 ;
        RECT 177.150 46.040 177.480 46.500 ;
        RECT 177.690 46.140 178.040 46.310 ;
        RECT 176.480 45.570 177.270 45.820 ;
        RECT 177.690 45.750 177.950 46.140 ;
        RECT 178.260 46.050 179.210 46.330 ;
        RECT 179.380 46.060 179.570 46.500 ;
        RECT 179.740 46.120 180.810 46.290 ;
        RECT 177.440 45.400 177.610 45.580 ;
        RECT 174.720 44.580 175.115 44.750 ;
        RECT 175.285 44.620 175.750 45.010 ;
        RECT 175.920 45.230 177.610 45.400 ;
        RECT 174.945 44.450 175.115 44.580 ;
        RECT 175.920 44.450 176.090 45.230 ;
        RECT 177.780 45.060 177.950 45.750 ;
        RECT 176.450 44.890 177.950 45.060 ;
        RECT 178.140 45.090 178.350 45.880 ;
        RECT 178.520 45.260 178.870 45.880 ;
        RECT 179.040 45.270 179.210 46.050 ;
        RECT 179.740 45.890 179.910 46.120 ;
        RECT 179.380 45.720 179.910 45.890 ;
        RECT 179.380 45.440 179.600 45.720 ;
        RECT 180.080 45.550 180.320 45.950 ;
        RECT 179.040 45.100 179.445 45.270 ;
        RECT 179.780 45.180 180.320 45.550 ;
        RECT 180.490 45.765 180.810 46.120 ;
        RECT 181.055 46.040 181.360 46.500 ;
        RECT 181.530 45.790 181.780 46.320 ;
        RECT 180.490 45.590 180.815 45.765 ;
        RECT 180.490 45.290 181.405 45.590 ;
        RECT 180.665 45.260 181.405 45.290 ;
        RECT 178.140 44.930 178.815 45.090 ;
        RECT 179.275 45.010 179.445 45.100 ;
        RECT 178.140 44.920 179.105 44.930 ;
        RECT 177.780 44.750 177.950 44.890 ;
        RECT 174.525 43.950 174.775 44.410 ;
        RECT 174.945 44.120 175.195 44.450 ;
        RECT 175.410 44.120 176.090 44.450 ;
        RECT 176.260 44.550 177.335 44.720 ;
        RECT 177.780 44.580 178.340 44.750 ;
        RECT 178.645 44.630 179.105 44.920 ;
        RECT 179.275 44.840 180.495 45.010 ;
        RECT 176.260 44.210 176.430 44.550 ;
        RECT 176.665 43.950 176.995 44.380 ;
        RECT 177.165 44.210 177.335 44.550 ;
        RECT 177.630 43.950 178.000 44.410 ;
        RECT 178.170 44.120 178.340 44.580 ;
        RECT 179.275 44.460 179.445 44.840 ;
        RECT 180.665 44.670 180.835 45.260 ;
        RECT 181.575 45.140 181.780 45.790 ;
        RECT 181.950 45.745 182.200 46.500 ;
        RECT 182.420 45.760 182.805 46.330 ;
        RECT 182.975 46.040 183.300 46.500 ;
        RECT 183.820 45.870 184.100 46.330 ;
        RECT 178.575 44.120 179.445 44.460 ;
        RECT 180.035 44.500 180.835 44.670 ;
        RECT 179.615 43.950 179.865 44.410 ;
        RECT 180.035 44.210 180.205 44.500 ;
        RECT 180.385 43.950 180.715 44.330 ;
        RECT 181.055 43.950 181.360 45.090 ;
        RECT 181.530 44.260 181.780 45.140 ;
        RECT 182.420 45.090 182.700 45.760 ;
        RECT 182.975 45.700 184.100 45.870 ;
        RECT 182.975 45.590 183.425 45.700 ;
        RECT 182.870 45.260 183.425 45.590 ;
        RECT 184.290 45.530 184.690 46.330 ;
        RECT 185.090 46.040 185.360 46.500 ;
        RECT 185.530 45.870 185.815 46.330 ;
        RECT 181.950 43.950 182.200 45.090 ;
        RECT 182.420 44.120 182.805 45.090 ;
        RECT 182.975 44.800 183.425 45.260 ;
        RECT 183.595 44.970 184.690 45.530 ;
        RECT 182.975 44.580 184.100 44.800 ;
        RECT 182.975 43.950 183.300 44.410 ;
        RECT 183.820 44.120 184.100 44.580 ;
        RECT 184.290 44.120 184.690 44.970 ;
        RECT 184.860 45.700 185.815 45.870 ;
        RECT 186.100 45.730 187.770 46.500 ;
        RECT 187.940 45.775 188.230 46.500 ;
        RECT 188.405 46.100 188.740 46.500 ;
        RECT 188.910 45.930 189.115 46.330 ;
        RECT 189.325 46.020 189.600 46.500 ;
        RECT 189.810 46.000 190.070 46.330 ;
        RECT 188.430 45.760 189.115 45.930 ;
        RECT 184.860 44.800 185.070 45.700 ;
        RECT 185.240 44.970 185.930 45.530 ;
        RECT 186.100 45.210 186.850 45.730 ;
        RECT 187.020 45.040 187.770 45.560 ;
        RECT 184.860 44.580 185.815 44.800 ;
        RECT 185.090 43.950 185.360 44.410 ;
        RECT 185.530 44.120 185.815 44.580 ;
        RECT 186.100 43.950 187.770 45.040 ;
        RECT 187.940 43.950 188.230 45.115 ;
        RECT 188.430 44.730 188.770 45.760 ;
        RECT 188.940 45.090 189.190 45.590 ;
        RECT 189.370 45.260 189.730 45.840 ;
        RECT 189.900 45.090 190.070 46.000 ;
        RECT 190.245 45.950 190.500 46.240 ;
        RECT 190.670 46.120 191.000 46.500 ;
        RECT 190.245 45.780 190.995 45.950 ;
        RECT 188.940 44.920 190.070 45.090 ;
        RECT 190.245 44.960 190.595 45.610 ;
        RECT 188.430 44.555 189.095 44.730 ;
        RECT 188.405 43.950 188.740 44.375 ;
        RECT 188.910 44.150 189.095 44.555 ;
        RECT 189.300 43.950 189.630 44.730 ;
        RECT 189.800 44.150 190.070 44.920 ;
        RECT 190.765 44.790 190.995 45.780 ;
        RECT 190.245 44.620 190.995 44.790 ;
        RECT 190.245 44.120 190.500 44.620 ;
        RECT 190.670 43.950 191.000 44.450 ;
        RECT 191.170 44.120 191.340 46.240 ;
        RECT 191.700 46.140 192.030 46.500 ;
        RECT 192.200 46.110 192.695 46.280 ;
        RECT 192.900 46.110 193.755 46.280 ;
        RECT 191.570 44.920 192.030 45.970 ;
        RECT 191.510 44.135 191.835 44.920 ;
        RECT 192.200 44.750 192.370 46.110 ;
        RECT 192.540 45.200 192.890 45.820 ;
        RECT 193.060 45.600 193.415 45.820 ;
        RECT 193.060 45.010 193.230 45.600 ;
        RECT 193.585 45.400 193.755 46.110 ;
        RECT 194.630 46.040 194.960 46.500 ;
        RECT 195.170 46.140 195.520 46.310 ;
        RECT 193.960 45.570 194.750 45.820 ;
        RECT 195.170 45.750 195.430 46.140 ;
        RECT 195.740 46.050 196.690 46.330 ;
        RECT 196.860 46.060 197.050 46.500 ;
        RECT 197.220 46.120 198.290 46.290 ;
        RECT 194.920 45.400 195.090 45.580 ;
        RECT 192.200 44.580 192.595 44.750 ;
        RECT 192.765 44.620 193.230 45.010 ;
        RECT 193.400 45.230 195.090 45.400 ;
        RECT 192.425 44.450 192.595 44.580 ;
        RECT 193.400 44.450 193.570 45.230 ;
        RECT 195.260 45.060 195.430 45.750 ;
        RECT 193.930 44.890 195.430 45.060 ;
        RECT 195.620 45.090 195.830 45.880 ;
        RECT 196.000 45.260 196.350 45.880 ;
        RECT 196.520 45.270 196.690 46.050 ;
        RECT 197.220 45.890 197.390 46.120 ;
        RECT 196.860 45.720 197.390 45.890 ;
        RECT 196.860 45.440 197.080 45.720 ;
        RECT 197.560 45.550 197.800 45.950 ;
        RECT 196.520 45.100 196.925 45.270 ;
        RECT 197.260 45.180 197.800 45.550 ;
        RECT 197.970 45.765 198.290 46.120 ;
        RECT 198.535 46.040 198.840 46.500 ;
        RECT 199.010 45.790 199.260 46.320 ;
        RECT 197.970 45.590 198.295 45.765 ;
        RECT 197.970 45.290 198.885 45.590 ;
        RECT 198.145 45.260 198.885 45.290 ;
        RECT 195.620 44.930 196.295 45.090 ;
        RECT 196.755 45.010 196.925 45.100 ;
        RECT 195.620 44.920 196.585 44.930 ;
        RECT 195.260 44.750 195.430 44.890 ;
        RECT 192.005 43.950 192.255 44.410 ;
        RECT 192.425 44.120 192.675 44.450 ;
        RECT 192.890 44.120 193.570 44.450 ;
        RECT 193.740 44.550 194.815 44.720 ;
        RECT 195.260 44.580 195.820 44.750 ;
        RECT 196.125 44.630 196.585 44.920 ;
        RECT 196.755 44.840 197.975 45.010 ;
        RECT 193.740 44.210 193.910 44.550 ;
        RECT 194.145 43.950 194.475 44.380 ;
        RECT 194.645 44.210 194.815 44.550 ;
        RECT 195.110 43.950 195.480 44.410 ;
        RECT 195.650 44.120 195.820 44.580 ;
        RECT 196.755 44.460 196.925 44.840 ;
        RECT 198.145 44.670 198.315 45.260 ;
        RECT 199.055 45.140 199.260 45.790 ;
        RECT 199.430 45.745 199.680 46.500 ;
        RECT 200.830 45.995 201.160 46.500 ;
        RECT 201.330 45.930 201.570 46.305 ;
        RECT 201.850 46.170 202.020 46.315 ;
        RECT 201.850 45.975 202.250 46.170 ;
        RECT 202.610 46.005 203.010 46.500 ;
        RECT 200.885 45.480 201.185 45.820 ;
        RECT 200.880 45.310 201.185 45.480 ;
        RECT 196.055 44.120 196.925 44.460 ;
        RECT 197.515 44.500 198.315 44.670 ;
        RECT 197.095 43.950 197.345 44.410 ;
        RECT 197.515 44.210 197.685 44.500 ;
        RECT 197.865 43.950 198.195 44.330 ;
        RECT 198.535 43.950 198.840 45.090 ;
        RECT 199.010 44.260 199.260 45.140 ;
        RECT 199.430 43.950 199.680 45.090 ;
        RECT 200.885 44.970 201.185 45.310 ;
        RECT 201.355 45.780 201.570 45.930 ;
        RECT 201.355 45.450 201.910 45.780 ;
        RECT 202.080 45.640 202.250 45.975 ;
        RECT 203.180 45.810 203.415 46.330 ;
        RECT 203.600 45.865 203.870 46.500 ;
        RECT 204.040 45.955 209.385 46.500 ;
        RECT 201.355 44.800 201.590 45.450 ;
        RECT 202.080 45.280 203.070 45.640 ;
        RECT 200.910 44.570 201.590 44.800 ;
        RECT 201.780 45.260 203.070 45.280 ;
        RECT 201.780 45.110 202.640 45.260 ;
        RECT 200.910 44.140 201.080 44.570 ;
        RECT 201.250 43.950 201.580 44.400 ;
        RECT 201.780 44.165 202.065 45.110 ;
        RECT 203.240 45.005 203.415 45.810 ;
        RECT 205.625 45.125 205.965 45.955 ;
        RECT 209.560 45.730 213.070 46.500 ;
        RECT 213.700 45.775 213.990 46.500 ;
        RECT 214.160 45.730 215.830 46.500 ;
        RECT 216.465 45.760 216.720 46.330 ;
        RECT 216.890 46.100 217.220 46.500 ;
        RECT 217.645 45.965 218.175 46.330 ;
        RECT 218.365 46.160 218.640 46.330 ;
        RECT 218.360 45.990 218.640 46.160 ;
        RECT 217.645 45.930 217.820 45.965 ;
        RECT 216.890 45.760 217.820 45.930 ;
        RECT 202.240 44.630 202.935 44.940 ;
        RECT 202.245 43.950 202.930 44.420 ;
        RECT 203.110 44.220 203.415 45.005 ;
        RECT 203.600 43.950 203.870 44.905 ;
        RECT 207.445 44.385 207.795 45.635 ;
        RECT 209.560 45.210 211.210 45.730 ;
        RECT 211.380 45.040 213.070 45.560 ;
        RECT 214.160 45.210 214.910 45.730 ;
        RECT 204.040 43.950 209.385 44.385 ;
        RECT 209.560 43.950 213.070 45.040 ;
        RECT 213.700 43.950 213.990 45.115 ;
        RECT 215.080 45.040 215.830 45.560 ;
        RECT 214.160 43.950 215.830 45.040 ;
        RECT 216.465 45.090 216.635 45.760 ;
        RECT 216.890 45.590 217.060 45.760 ;
        RECT 216.805 45.260 217.060 45.590 ;
        RECT 217.285 45.260 217.480 45.590 ;
        RECT 216.465 44.120 216.800 45.090 ;
        RECT 216.970 43.950 217.140 45.090 ;
        RECT 217.310 44.290 217.480 45.260 ;
        RECT 217.650 44.630 217.820 45.760 ;
        RECT 217.990 44.970 218.160 45.770 ;
        RECT 218.365 45.170 218.640 45.990 ;
        RECT 218.810 44.970 219.000 46.330 ;
        RECT 219.180 45.965 219.690 46.500 ;
        RECT 219.910 45.690 220.155 46.295 ;
        RECT 222.040 46.030 222.340 46.500 ;
        RECT 222.510 45.860 222.765 46.305 ;
        RECT 222.935 46.030 223.195 46.500 ;
        RECT 223.365 45.860 223.625 46.305 ;
        RECT 223.795 46.030 224.090 46.500 ;
        RECT 221.520 45.690 224.550 45.860 ;
        RECT 219.200 45.520 220.430 45.690 ;
        RECT 217.990 44.800 219.000 44.970 ;
        RECT 219.170 44.955 219.920 45.145 ;
        RECT 217.650 44.460 218.775 44.630 ;
        RECT 219.170 44.290 219.340 44.955 ;
        RECT 220.090 44.710 220.430 45.520 ;
        RECT 221.520 45.125 221.820 45.690 ;
        RECT 221.995 45.295 224.210 45.520 ;
        RECT 224.380 45.125 224.550 45.690 ;
        RECT 221.520 44.955 224.550 45.125 ;
        RECT 224.740 45.760 225.125 46.330 ;
        RECT 225.295 46.040 225.620 46.500 ;
        RECT 226.140 45.870 226.420 46.330 ;
        RECT 224.740 45.090 225.020 45.760 ;
        RECT 225.295 45.700 226.420 45.870 ;
        RECT 225.295 45.590 225.745 45.700 ;
        RECT 225.190 45.260 225.745 45.590 ;
        RECT 226.610 45.530 227.010 46.330 ;
        RECT 227.410 46.040 227.680 46.500 ;
        RECT 227.850 45.870 228.135 46.330 ;
        RECT 217.310 44.120 219.340 44.290 ;
        RECT 219.510 43.950 219.680 44.710 ;
        RECT 219.915 44.300 220.430 44.710 ;
        RECT 221.520 43.950 221.905 44.785 ;
        RECT 222.075 44.150 222.335 44.955 ;
        RECT 222.505 43.950 222.765 44.785 ;
        RECT 222.935 44.150 223.190 44.955 ;
        RECT 223.365 43.950 223.625 44.785 ;
        RECT 223.795 44.150 224.050 44.955 ;
        RECT 224.225 43.950 224.570 44.785 ;
        RECT 224.740 44.120 225.125 45.090 ;
        RECT 225.295 44.800 225.745 45.260 ;
        RECT 225.915 44.970 227.010 45.530 ;
        RECT 225.295 44.580 226.420 44.800 ;
        RECT 225.295 43.950 225.620 44.410 ;
        RECT 226.140 44.120 226.420 44.580 ;
        RECT 226.610 44.120 227.010 44.970 ;
        RECT 227.180 45.700 228.135 45.870 ;
        RECT 228.510 45.950 228.680 46.330 ;
        RECT 228.895 46.120 229.225 46.500 ;
        RECT 228.510 45.780 229.225 45.950 ;
        RECT 227.180 44.800 227.390 45.700 ;
        RECT 227.560 44.970 228.250 45.530 ;
        RECT 228.420 45.230 228.775 45.600 ;
        RECT 229.055 45.590 229.225 45.780 ;
        RECT 229.395 45.755 229.650 46.330 ;
        RECT 229.055 45.260 229.310 45.590 ;
        RECT 229.055 45.050 229.225 45.260 ;
        RECT 228.510 44.880 229.225 45.050 ;
        RECT 229.480 45.025 229.650 45.755 ;
        RECT 229.825 45.660 230.085 46.500 ;
        RECT 230.265 45.950 230.520 46.240 ;
        RECT 230.690 46.120 231.020 46.500 ;
        RECT 230.265 45.780 231.015 45.950 ;
        RECT 227.180 44.580 228.135 44.800 ;
        RECT 227.410 43.950 227.680 44.410 ;
        RECT 227.850 44.120 228.135 44.580 ;
        RECT 228.510 44.120 228.680 44.880 ;
        RECT 228.895 43.950 229.225 44.710 ;
        RECT 229.395 44.120 229.650 45.025 ;
        RECT 229.825 43.950 230.085 45.100 ;
        RECT 230.265 44.960 230.615 45.610 ;
        RECT 230.785 44.790 231.015 45.780 ;
        RECT 230.265 44.620 231.015 44.790 ;
        RECT 230.265 44.120 230.520 44.620 ;
        RECT 230.690 43.950 231.020 44.450 ;
        RECT 231.190 44.120 231.360 46.240 ;
        RECT 231.720 46.140 232.050 46.500 ;
        RECT 232.220 46.110 232.715 46.280 ;
        RECT 232.920 46.110 233.775 46.280 ;
        RECT 231.590 44.920 232.050 45.970 ;
        RECT 231.530 44.135 231.855 44.920 ;
        RECT 232.220 44.750 232.390 46.110 ;
        RECT 232.560 45.200 232.910 45.820 ;
        RECT 233.080 45.600 233.435 45.820 ;
        RECT 233.080 45.010 233.250 45.600 ;
        RECT 233.605 45.400 233.775 46.110 ;
        RECT 234.650 46.040 234.980 46.500 ;
        RECT 235.190 46.140 235.540 46.310 ;
        RECT 233.980 45.570 234.770 45.820 ;
        RECT 235.190 45.750 235.450 46.140 ;
        RECT 235.760 46.050 236.710 46.330 ;
        RECT 236.880 46.060 237.070 46.500 ;
        RECT 237.240 46.120 238.310 46.290 ;
        RECT 234.940 45.400 235.110 45.580 ;
        RECT 232.220 44.580 232.615 44.750 ;
        RECT 232.785 44.620 233.250 45.010 ;
        RECT 233.420 45.230 235.110 45.400 ;
        RECT 232.445 44.450 232.615 44.580 ;
        RECT 233.420 44.450 233.590 45.230 ;
        RECT 235.280 45.060 235.450 45.750 ;
        RECT 233.950 44.890 235.450 45.060 ;
        RECT 235.640 45.090 235.850 45.880 ;
        RECT 236.020 45.260 236.370 45.880 ;
        RECT 236.540 45.270 236.710 46.050 ;
        RECT 237.240 45.890 237.410 46.120 ;
        RECT 236.880 45.720 237.410 45.890 ;
        RECT 236.880 45.440 237.100 45.720 ;
        RECT 237.580 45.550 237.820 45.950 ;
        RECT 236.540 45.100 236.945 45.270 ;
        RECT 237.280 45.180 237.820 45.550 ;
        RECT 237.990 45.765 238.310 46.120 ;
        RECT 238.555 46.040 238.860 46.500 ;
        RECT 239.030 45.790 239.285 46.320 ;
        RECT 237.990 45.590 238.315 45.765 ;
        RECT 237.990 45.290 238.905 45.590 ;
        RECT 238.165 45.260 238.905 45.290 ;
        RECT 235.640 44.930 236.315 45.090 ;
        RECT 236.775 45.010 236.945 45.100 ;
        RECT 235.640 44.920 236.605 44.930 ;
        RECT 235.280 44.750 235.450 44.890 ;
        RECT 232.025 43.950 232.275 44.410 ;
        RECT 232.445 44.120 232.695 44.450 ;
        RECT 232.910 44.120 233.590 44.450 ;
        RECT 233.760 44.550 234.835 44.720 ;
        RECT 235.280 44.580 235.840 44.750 ;
        RECT 236.145 44.630 236.605 44.920 ;
        RECT 236.775 44.840 237.995 45.010 ;
        RECT 233.760 44.210 233.930 44.550 ;
        RECT 234.165 43.950 234.495 44.380 ;
        RECT 234.665 44.210 234.835 44.550 ;
        RECT 235.130 43.950 235.500 44.410 ;
        RECT 235.670 44.120 235.840 44.580 ;
        RECT 236.775 44.460 236.945 44.840 ;
        RECT 238.165 44.670 238.335 45.260 ;
        RECT 239.075 45.140 239.285 45.790 ;
        RECT 239.460 45.775 239.750 46.500 ;
        RECT 236.075 44.120 236.945 44.460 ;
        RECT 237.535 44.500 238.335 44.670 ;
        RECT 237.115 43.950 237.365 44.410 ;
        RECT 237.535 44.210 237.705 44.500 ;
        RECT 237.885 43.950 238.215 44.330 ;
        RECT 238.555 43.950 238.860 45.090 ;
        RECT 239.030 44.260 239.285 45.140 ;
        RECT 239.920 45.680 240.605 46.320 ;
        RECT 240.775 45.680 240.945 46.500 ;
        RECT 241.115 45.850 241.445 46.315 ;
        RECT 241.615 46.030 241.785 46.500 ;
        RECT 242.045 46.110 243.230 46.280 ;
        RECT 243.400 45.940 243.730 46.330 ;
        RECT 242.430 45.850 242.815 45.940 ;
        RECT 241.115 45.680 242.815 45.850 ;
        RECT 243.220 45.760 243.730 45.940 ;
        RECT 244.060 45.760 244.445 46.330 ;
        RECT 244.615 46.040 244.940 46.500 ;
        RECT 245.460 45.870 245.740 46.330 ;
        RECT 239.460 43.950 239.750 45.115 ;
        RECT 239.920 44.710 240.170 45.680 ;
        RECT 240.340 45.300 240.675 45.510 ;
        RECT 240.845 45.300 241.295 45.510 ;
        RECT 241.485 45.480 241.970 45.510 ;
        RECT 241.485 45.310 241.990 45.480 ;
        RECT 241.485 45.300 241.970 45.310 ;
        RECT 240.505 45.130 240.675 45.300 ;
        RECT 240.505 44.960 241.425 45.130 ;
        RECT 239.920 44.120 240.585 44.710 ;
        RECT 240.755 43.950 241.085 44.790 ;
        RECT 241.255 44.710 241.425 44.960 ;
        RECT 241.595 44.880 241.970 45.300 ;
        RECT 242.160 45.260 242.540 45.510 ;
        RECT 242.720 45.300 243.050 45.510 ;
        RECT 242.160 44.880 242.480 45.260 ;
        RECT 243.220 45.130 243.390 45.760 ;
        RECT 243.560 45.300 243.890 45.590 ;
        RECT 242.650 44.960 243.735 45.130 ;
        RECT 242.650 44.710 242.820 44.960 ;
        RECT 241.255 44.540 242.820 44.710 ;
        RECT 241.595 44.120 242.400 44.540 ;
        RECT 242.990 43.950 243.240 44.790 ;
        RECT 243.435 44.120 243.735 44.960 ;
        RECT 244.060 45.090 244.340 45.760 ;
        RECT 244.615 45.700 245.740 45.870 ;
        RECT 244.615 45.590 245.065 45.700 ;
        RECT 244.510 45.260 245.065 45.590 ;
        RECT 245.930 45.530 246.330 46.330 ;
        RECT 246.730 46.040 247.000 46.500 ;
        RECT 247.170 45.870 247.455 46.330 ;
        RECT 244.060 44.120 244.445 45.090 ;
        RECT 244.615 44.800 245.065 45.260 ;
        RECT 245.235 44.970 246.330 45.530 ;
        RECT 244.615 44.580 245.740 44.800 ;
        RECT 244.615 43.950 244.940 44.410 ;
        RECT 245.460 44.120 245.740 44.580 ;
        RECT 245.930 44.120 246.330 44.970 ;
        RECT 246.500 45.700 247.455 45.870 ;
        RECT 248.205 45.950 248.460 46.240 ;
        RECT 248.630 46.120 248.960 46.500 ;
        RECT 248.205 45.780 248.955 45.950 ;
        RECT 246.500 44.800 246.710 45.700 ;
        RECT 246.880 44.970 247.570 45.530 ;
        RECT 248.205 44.960 248.555 45.610 ;
        RECT 246.500 44.580 247.455 44.800 ;
        RECT 248.725 44.790 248.955 45.780 ;
        RECT 246.730 43.950 247.000 44.410 ;
        RECT 247.170 44.120 247.455 44.580 ;
        RECT 248.205 44.620 248.955 44.790 ;
        RECT 248.205 44.120 248.460 44.620 ;
        RECT 248.630 43.950 248.960 44.450 ;
        RECT 249.130 44.120 249.300 46.240 ;
        RECT 249.660 46.140 249.990 46.500 ;
        RECT 250.160 46.110 250.655 46.280 ;
        RECT 250.860 46.110 251.715 46.280 ;
        RECT 249.530 44.920 249.990 45.970 ;
        RECT 249.470 44.135 249.795 44.920 ;
        RECT 250.160 44.750 250.330 46.110 ;
        RECT 250.500 45.200 250.850 45.820 ;
        RECT 251.020 45.600 251.375 45.820 ;
        RECT 251.020 45.010 251.190 45.600 ;
        RECT 251.545 45.400 251.715 46.110 ;
        RECT 252.590 46.040 252.920 46.500 ;
        RECT 253.130 46.140 253.480 46.310 ;
        RECT 251.920 45.570 252.710 45.820 ;
        RECT 253.130 45.750 253.390 46.140 ;
        RECT 253.700 46.050 254.650 46.330 ;
        RECT 254.820 46.060 255.010 46.500 ;
        RECT 255.180 46.120 256.250 46.290 ;
        RECT 252.880 45.400 253.050 45.580 ;
        RECT 250.160 44.580 250.555 44.750 ;
        RECT 250.725 44.620 251.190 45.010 ;
        RECT 251.360 45.230 253.050 45.400 ;
        RECT 250.385 44.450 250.555 44.580 ;
        RECT 251.360 44.450 251.530 45.230 ;
        RECT 253.220 45.060 253.390 45.750 ;
        RECT 251.890 44.890 253.390 45.060 ;
        RECT 253.580 45.090 253.790 45.880 ;
        RECT 253.960 45.260 254.310 45.880 ;
        RECT 254.480 45.270 254.650 46.050 ;
        RECT 255.180 45.890 255.350 46.120 ;
        RECT 254.820 45.720 255.350 45.890 ;
        RECT 254.820 45.440 255.040 45.720 ;
        RECT 255.520 45.550 255.760 45.950 ;
        RECT 254.480 45.100 254.885 45.270 ;
        RECT 255.220 45.180 255.760 45.550 ;
        RECT 255.930 45.765 256.250 46.120 ;
        RECT 256.495 46.040 256.800 46.500 ;
        RECT 256.970 45.790 257.225 46.320 ;
        RECT 255.930 45.590 256.255 45.765 ;
        RECT 255.930 45.290 256.845 45.590 ;
        RECT 256.105 45.260 256.845 45.290 ;
        RECT 253.580 44.930 254.255 45.090 ;
        RECT 254.715 45.010 254.885 45.100 ;
        RECT 253.580 44.920 254.545 44.930 ;
        RECT 253.220 44.750 253.390 44.890 ;
        RECT 249.965 43.950 250.215 44.410 ;
        RECT 250.385 44.120 250.635 44.450 ;
        RECT 250.850 44.120 251.530 44.450 ;
        RECT 251.700 44.550 252.775 44.720 ;
        RECT 253.220 44.580 253.780 44.750 ;
        RECT 254.085 44.630 254.545 44.920 ;
        RECT 254.715 44.840 255.935 45.010 ;
        RECT 251.700 44.210 251.870 44.550 ;
        RECT 252.105 43.950 252.435 44.380 ;
        RECT 252.605 44.210 252.775 44.550 ;
        RECT 253.070 43.950 253.440 44.410 ;
        RECT 253.610 44.120 253.780 44.580 ;
        RECT 254.715 44.460 254.885 44.840 ;
        RECT 256.105 44.670 256.275 45.260 ;
        RECT 257.015 45.140 257.225 45.790 ;
        RECT 254.015 44.120 254.885 44.460 ;
        RECT 255.475 44.500 256.275 44.670 ;
        RECT 255.055 43.950 255.305 44.410 ;
        RECT 255.475 44.210 255.645 44.500 ;
        RECT 255.825 43.950 256.155 44.330 ;
        RECT 256.495 43.950 256.800 45.090 ;
        RECT 256.970 44.260 257.225 45.140 ;
        RECT 257.400 45.680 258.085 46.320 ;
        RECT 258.255 45.680 258.425 46.500 ;
        RECT 258.595 45.850 258.925 46.315 ;
        RECT 259.095 46.030 259.265 46.500 ;
        RECT 259.525 46.110 260.710 46.280 ;
        RECT 260.880 45.940 261.210 46.330 ;
        RECT 259.910 45.850 260.295 45.940 ;
        RECT 258.595 45.680 260.295 45.850 ;
        RECT 260.700 45.760 261.210 45.940 ;
        RECT 261.540 45.760 261.925 46.330 ;
        RECT 262.095 46.040 262.420 46.500 ;
        RECT 262.940 45.870 263.220 46.330 ;
        RECT 257.400 44.710 257.650 45.680 ;
        RECT 257.820 45.300 258.155 45.510 ;
        RECT 258.325 45.300 258.775 45.510 ;
        RECT 258.965 45.480 259.450 45.510 ;
        RECT 258.965 45.310 259.470 45.480 ;
        RECT 258.965 45.300 259.450 45.310 ;
        RECT 257.985 45.130 258.155 45.300 ;
        RECT 257.985 44.960 258.905 45.130 ;
        RECT 257.400 44.120 258.065 44.710 ;
        RECT 258.235 43.950 258.565 44.790 ;
        RECT 258.735 44.710 258.905 44.960 ;
        RECT 259.075 44.880 259.450 45.300 ;
        RECT 259.640 45.260 260.020 45.510 ;
        RECT 260.200 45.300 260.530 45.510 ;
        RECT 259.640 44.880 259.960 45.260 ;
        RECT 260.700 45.130 260.870 45.760 ;
        RECT 261.040 45.300 261.370 45.590 ;
        RECT 260.130 44.960 261.215 45.130 ;
        RECT 260.130 44.710 260.300 44.960 ;
        RECT 258.735 44.540 260.300 44.710 ;
        RECT 259.075 44.120 259.880 44.540 ;
        RECT 260.470 43.950 260.720 44.790 ;
        RECT 260.915 44.120 261.215 44.960 ;
        RECT 261.540 45.090 261.820 45.760 ;
        RECT 262.095 45.700 263.220 45.870 ;
        RECT 262.095 45.590 262.545 45.700 ;
        RECT 261.990 45.260 262.545 45.590 ;
        RECT 263.410 45.530 263.810 46.330 ;
        RECT 264.210 46.040 264.480 46.500 ;
        RECT 264.650 45.870 264.935 46.330 ;
        RECT 261.540 44.120 261.925 45.090 ;
        RECT 262.095 44.800 262.545 45.260 ;
        RECT 262.715 44.970 263.810 45.530 ;
        RECT 262.095 44.580 263.220 44.800 ;
        RECT 262.095 43.950 262.420 44.410 ;
        RECT 262.940 44.120 263.220 44.580 ;
        RECT 263.410 44.120 263.810 44.970 ;
        RECT 263.980 45.700 264.935 45.870 ;
        RECT 265.220 45.775 265.510 46.500 ;
        RECT 265.715 45.760 266.330 46.330 ;
        RECT 266.500 45.990 266.715 46.500 ;
        RECT 266.945 45.990 267.225 46.320 ;
        RECT 267.405 45.990 267.645 46.500 ;
        RECT 263.980 44.800 264.190 45.700 ;
        RECT 264.360 44.970 265.050 45.530 ;
        RECT 263.980 44.580 264.935 44.800 ;
        RECT 264.210 43.950 264.480 44.410 ;
        RECT 264.650 44.120 264.935 44.580 ;
        RECT 265.220 43.950 265.510 45.115 ;
        RECT 265.715 44.740 266.030 45.760 ;
        RECT 266.200 45.090 266.370 45.590 ;
        RECT 266.620 45.260 266.885 45.820 ;
        RECT 267.055 45.090 267.225 45.990 ;
        RECT 267.395 45.260 267.750 45.820 ;
        RECT 268.020 45.680 268.250 46.500 ;
        RECT 268.420 45.700 268.750 46.330 ;
        RECT 268.000 45.260 268.330 45.510 ;
        RECT 268.500 45.100 268.750 45.700 ;
        RECT 268.920 45.680 269.130 46.500 ;
        RECT 269.360 45.730 271.030 46.500 ;
        RECT 271.665 45.970 271.955 46.320 ;
        RECT 272.150 46.140 272.480 46.500 ;
        RECT 272.650 45.970 272.880 46.275 ;
        RECT 271.665 45.800 272.880 45.970 ;
        RECT 273.070 46.160 273.240 46.195 ;
        RECT 273.070 45.990 273.270 46.160 ;
        RECT 269.360 45.210 270.110 45.730 ;
        RECT 273.070 45.630 273.240 45.990 ;
        RECT 266.200 44.920 267.625 45.090 ;
        RECT 265.715 44.120 266.250 44.740 ;
        RECT 266.420 43.950 266.750 44.750 ;
        RECT 267.235 44.745 267.625 44.920 ;
        RECT 268.020 43.950 268.250 45.090 ;
        RECT 268.420 44.120 268.750 45.100 ;
        RECT 268.920 43.950 269.130 45.090 ;
        RECT 270.280 45.040 271.030 45.560 ;
        RECT 271.725 45.480 271.985 45.590 ;
        RECT 271.720 45.310 271.985 45.480 ;
        RECT 271.725 45.260 271.985 45.310 ;
        RECT 272.165 45.260 272.550 45.590 ;
        RECT 272.720 45.460 273.240 45.630 ;
        RECT 273.960 45.760 274.345 46.330 ;
        RECT 274.515 46.040 274.840 46.500 ;
        RECT 275.360 45.870 275.640 46.330 ;
        RECT 269.360 43.950 271.030 45.040 ;
        RECT 271.665 43.950 271.985 45.090 ;
        RECT 272.165 44.210 272.360 45.260 ;
        RECT 272.720 45.080 272.890 45.460 ;
        RECT 272.540 44.800 272.890 45.080 ;
        RECT 273.080 44.930 273.325 45.290 ;
        RECT 273.960 45.090 274.240 45.760 ;
        RECT 274.515 45.700 275.640 45.870 ;
        RECT 274.515 45.590 274.965 45.700 ;
        RECT 274.410 45.260 274.965 45.590 ;
        RECT 275.830 45.530 276.230 46.330 ;
        RECT 276.630 46.040 276.900 46.500 ;
        RECT 277.070 45.870 277.355 46.330 ;
        RECT 272.540 44.120 272.870 44.800 ;
        RECT 273.070 43.950 273.325 44.750 ;
        RECT 273.960 44.120 274.345 45.090 ;
        RECT 274.515 44.800 274.965 45.260 ;
        RECT 275.135 44.970 276.230 45.530 ;
        RECT 274.515 44.580 275.640 44.800 ;
        RECT 274.515 43.950 274.840 44.410 ;
        RECT 275.360 44.120 275.640 44.580 ;
        RECT 275.830 44.120 276.230 44.970 ;
        RECT 276.400 45.700 277.355 45.870 ;
        RECT 277.640 45.750 278.850 46.500 ;
        RECT 279.135 45.870 279.420 46.330 ;
        RECT 279.590 46.040 279.860 46.500 ;
        RECT 276.400 44.800 276.610 45.700 ;
        RECT 276.780 44.970 277.470 45.530 ;
        RECT 277.640 45.210 278.160 45.750 ;
        RECT 279.135 45.700 280.090 45.870 ;
        RECT 278.330 45.040 278.850 45.580 ;
        RECT 276.400 44.580 277.355 44.800 ;
        RECT 276.630 43.950 276.900 44.410 ;
        RECT 277.070 44.120 277.355 44.580 ;
        RECT 277.640 43.950 278.850 45.040 ;
        RECT 279.020 44.970 279.710 45.530 ;
        RECT 279.880 44.800 280.090 45.700 ;
        RECT 279.135 44.580 280.090 44.800 ;
        RECT 280.260 45.530 280.660 46.330 ;
        RECT 280.850 45.870 281.130 46.330 ;
        RECT 281.650 46.040 281.975 46.500 ;
        RECT 280.850 45.700 281.975 45.870 ;
        RECT 282.145 45.760 282.530 46.330 ;
        RECT 282.700 45.955 288.045 46.500 ;
        RECT 281.525 45.590 281.975 45.700 ;
        RECT 280.260 44.970 281.355 45.530 ;
        RECT 281.525 45.260 282.080 45.590 ;
        RECT 279.135 44.120 279.420 44.580 ;
        RECT 279.590 43.950 279.860 44.410 ;
        RECT 280.260 44.120 280.660 44.970 ;
        RECT 281.525 44.800 281.975 45.260 ;
        RECT 282.250 45.090 282.530 45.760 ;
        RECT 284.285 45.125 284.625 45.955 ;
        RECT 288.220 45.730 290.810 46.500 ;
        RECT 290.980 45.775 291.270 46.500 ;
        RECT 291.440 45.730 294.950 46.500 ;
        RECT 295.120 45.750 296.330 46.500 ;
        RECT 296.505 45.950 296.760 46.240 ;
        RECT 296.930 46.120 297.260 46.500 ;
        RECT 296.505 45.780 297.255 45.950 ;
        RECT 280.850 44.580 281.975 44.800 ;
        RECT 280.850 44.120 281.130 44.580 ;
        RECT 281.650 43.950 281.975 44.410 ;
        RECT 282.145 44.120 282.530 45.090 ;
        RECT 286.105 44.385 286.455 45.635 ;
        RECT 288.220 45.210 289.430 45.730 ;
        RECT 289.600 45.040 290.810 45.560 ;
        RECT 291.440 45.210 293.090 45.730 ;
        RECT 282.700 43.950 288.045 44.385 ;
        RECT 288.220 43.950 290.810 45.040 ;
        RECT 290.980 43.950 291.270 45.115 ;
        RECT 293.260 45.040 294.950 45.560 ;
        RECT 295.120 45.210 295.640 45.750 ;
        RECT 295.810 45.040 296.330 45.580 ;
        RECT 291.440 43.950 294.950 45.040 ;
        RECT 295.120 43.950 296.330 45.040 ;
        RECT 296.505 44.960 296.855 45.610 ;
        RECT 297.025 44.790 297.255 45.780 ;
        RECT 296.505 44.620 297.255 44.790 ;
        RECT 296.505 44.120 296.760 44.620 ;
        RECT 296.930 43.950 297.260 44.450 ;
        RECT 297.430 44.120 297.600 46.240 ;
        RECT 297.960 46.140 298.290 46.500 ;
        RECT 298.460 46.110 298.955 46.280 ;
        RECT 299.160 46.110 300.015 46.280 ;
        RECT 297.830 44.920 298.290 45.970 ;
        RECT 297.770 44.135 298.095 44.920 ;
        RECT 298.460 44.750 298.630 46.110 ;
        RECT 298.800 45.200 299.150 45.820 ;
        RECT 299.320 45.600 299.675 45.820 ;
        RECT 299.320 45.010 299.490 45.600 ;
        RECT 299.845 45.400 300.015 46.110 ;
        RECT 300.890 46.040 301.220 46.500 ;
        RECT 301.430 46.140 301.780 46.310 ;
        RECT 300.220 45.570 301.010 45.820 ;
        RECT 301.430 45.750 301.690 46.140 ;
        RECT 302.000 46.050 302.950 46.330 ;
        RECT 303.120 46.060 303.310 46.500 ;
        RECT 303.480 46.120 304.550 46.290 ;
        RECT 301.180 45.400 301.350 45.580 ;
        RECT 298.460 44.580 298.855 44.750 ;
        RECT 299.025 44.620 299.490 45.010 ;
        RECT 299.660 45.230 301.350 45.400 ;
        RECT 298.685 44.450 298.855 44.580 ;
        RECT 299.660 44.450 299.830 45.230 ;
        RECT 301.520 45.060 301.690 45.750 ;
        RECT 300.190 44.890 301.690 45.060 ;
        RECT 301.880 45.090 302.090 45.880 ;
        RECT 302.260 45.260 302.610 45.880 ;
        RECT 302.780 45.270 302.950 46.050 ;
        RECT 303.480 45.890 303.650 46.120 ;
        RECT 303.120 45.720 303.650 45.890 ;
        RECT 303.120 45.440 303.340 45.720 ;
        RECT 303.820 45.550 304.060 45.950 ;
        RECT 302.780 45.100 303.185 45.270 ;
        RECT 303.520 45.180 304.060 45.550 ;
        RECT 304.230 45.765 304.550 46.120 ;
        RECT 304.795 46.040 305.100 46.500 ;
        RECT 305.270 45.790 305.525 46.320 ;
        RECT 304.230 45.590 304.555 45.765 ;
        RECT 304.230 45.290 305.145 45.590 ;
        RECT 304.405 45.260 305.145 45.290 ;
        RECT 301.880 44.930 302.555 45.090 ;
        RECT 303.015 45.010 303.185 45.100 ;
        RECT 301.880 44.920 302.845 44.930 ;
        RECT 301.520 44.750 301.690 44.890 ;
        RECT 298.265 43.950 298.515 44.410 ;
        RECT 298.685 44.120 298.935 44.450 ;
        RECT 299.150 44.120 299.830 44.450 ;
        RECT 300.000 44.550 301.075 44.720 ;
        RECT 301.520 44.580 302.080 44.750 ;
        RECT 302.385 44.630 302.845 44.920 ;
        RECT 303.015 44.840 304.235 45.010 ;
        RECT 300.000 44.210 300.170 44.550 ;
        RECT 300.405 43.950 300.735 44.380 ;
        RECT 300.905 44.210 301.075 44.550 ;
        RECT 301.370 43.950 301.740 44.410 ;
        RECT 301.910 44.120 302.080 44.580 ;
        RECT 303.015 44.460 303.185 44.840 ;
        RECT 304.405 44.670 304.575 45.260 ;
        RECT 305.315 45.140 305.525 45.790 ;
        RECT 305.700 45.730 307.370 46.500 ;
        RECT 308.090 45.950 308.260 46.330 ;
        RECT 308.475 46.120 308.805 46.500 ;
        RECT 308.090 45.780 308.805 45.950 ;
        RECT 305.700 45.210 306.450 45.730 ;
        RECT 302.315 44.120 303.185 44.460 ;
        RECT 303.775 44.500 304.575 44.670 ;
        RECT 303.355 43.950 303.605 44.410 ;
        RECT 303.775 44.210 303.945 44.500 ;
        RECT 304.125 43.950 304.455 44.330 ;
        RECT 304.795 43.950 305.100 45.090 ;
        RECT 305.270 44.260 305.525 45.140 ;
        RECT 306.620 45.040 307.370 45.560 ;
        RECT 308.000 45.230 308.355 45.600 ;
        RECT 308.635 45.590 308.805 45.780 ;
        RECT 308.975 45.755 309.230 46.330 ;
        RECT 308.635 45.260 308.890 45.590 ;
        RECT 308.635 45.050 308.805 45.260 ;
        RECT 305.700 43.950 307.370 45.040 ;
        RECT 308.090 44.880 308.805 45.050 ;
        RECT 309.060 45.025 309.230 45.755 ;
        RECT 309.405 45.660 309.665 46.500 ;
        RECT 309.840 45.750 311.050 46.500 ;
        RECT 308.090 44.120 308.260 44.880 ;
        RECT 308.475 43.950 308.805 44.710 ;
        RECT 308.975 44.120 309.230 45.025 ;
        RECT 309.405 43.950 309.665 45.100 ;
        RECT 309.840 45.040 310.360 45.580 ;
        RECT 310.530 45.210 311.050 45.750 ;
        RECT 309.840 43.950 311.050 45.040 ;
        RECT 162.095 43.780 311.135 43.950 ;
        RECT 162.180 42.690 163.390 43.780 ;
        RECT 163.560 42.690 165.230 43.780 ;
        RECT 165.865 43.110 166.120 43.610 ;
        RECT 166.290 43.280 166.620 43.780 ;
        RECT 165.865 42.940 166.615 43.110 ;
        RECT 162.180 41.980 162.700 42.520 ;
        RECT 162.870 42.150 163.390 42.690 ;
        RECT 163.560 42.000 164.310 42.520 ;
        RECT 164.480 42.170 165.230 42.690 ;
        RECT 165.865 42.120 166.215 42.770 ;
        RECT 162.180 41.230 163.390 41.980 ;
        RECT 163.560 41.230 165.230 42.000 ;
        RECT 166.385 41.950 166.615 42.940 ;
        RECT 165.865 41.780 166.615 41.950 ;
        RECT 165.865 41.490 166.120 41.780 ;
        RECT 166.290 41.230 166.620 41.610 ;
        RECT 166.790 41.490 166.960 43.610 ;
        RECT 167.130 42.810 167.455 43.595 ;
        RECT 167.625 43.320 167.875 43.780 ;
        RECT 168.045 43.280 168.295 43.610 ;
        RECT 168.510 43.280 169.190 43.610 ;
        RECT 168.045 43.150 168.215 43.280 ;
        RECT 167.820 42.980 168.215 43.150 ;
        RECT 167.190 41.760 167.650 42.810 ;
        RECT 167.820 41.620 167.990 42.980 ;
        RECT 168.385 42.720 168.850 43.110 ;
        RECT 168.160 41.910 168.510 42.530 ;
        RECT 168.680 42.130 168.850 42.720 ;
        RECT 169.020 42.500 169.190 43.280 ;
        RECT 169.360 43.180 169.530 43.520 ;
        RECT 169.765 43.350 170.095 43.780 ;
        RECT 170.265 43.180 170.435 43.520 ;
        RECT 170.730 43.320 171.100 43.780 ;
        RECT 169.360 43.010 170.435 43.180 ;
        RECT 171.270 43.150 171.440 43.610 ;
        RECT 171.675 43.270 172.545 43.610 ;
        RECT 172.715 43.320 172.965 43.780 ;
        RECT 170.880 42.980 171.440 43.150 ;
        RECT 170.880 42.840 171.050 42.980 ;
        RECT 169.550 42.670 171.050 42.840 ;
        RECT 171.745 42.810 172.205 43.100 ;
        RECT 169.020 42.330 170.710 42.500 ;
        RECT 168.680 41.910 169.035 42.130 ;
        RECT 169.205 41.620 169.375 42.330 ;
        RECT 169.580 41.910 170.370 42.160 ;
        RECT 170.540 42.150 170.710 42.330 ;
        RECT 170.880 41.980 171.050 42.670 ;
        RECT 167.320 41.230 167.650 41.590 ;
        RECT 167.820 41.450 168.315 41.620 ;
        RECT 168.520 41.450 169.375 41.620 ;
        RECT 170.250 41.230 170.580 41.690 ;
        RECT 170.790 41.590 171.050 41.980 ;
        RECT 171.240 42.800 172.205 42.810 ;
        RECT 172.375 42.890 172.545 43.270 ;
        RECT 173.135 43.230 173.305 43.520 ;
        RECT 173.485 43.400 173.815 43.780 ;
        RECT 173.135 43.060 173.935 43.230 ;
        RECT 171.240 42.640 171.915 42.800 ;
        RECT 172.375 42.720 173.595 42.890 ;
        RECT 171.240 41.850 171.450 42.640 ;
        RECT 172.375 42.630 172.545 42.720 ;
        RECT 171.620 41.850 171.970 42.470 ;
        RECT 172.140 42.460 172.545 42.630 ;
        RECT 172.140 41.680 172.310 42.460 ;
        RECT 172.480 42.010 172.700 42.290 ;
        RECT 172.880 42.180 173.420 42.550 ;
        RECT 173.765 42.470 173.935 43.060 ;
        RECT 174.155 42.640 174.460 43.780 ;
        RECT 174.630 42.590 174.885 43.470 ;
        RECT 175.060 42.615 175.350 43.780 ;
        RECT 175.525 43.110 175.780 43.610 ;
        RECT 175.950 43.280 176.280 43.780 ;
        RECT 175.525 42.940 176.275 43.110 ;
        RECT 173.765 42.440 174.505 42.470 ;
        RECT 172.480 41.840 173.010 42.010 ;
        RECT 170.790 41.420 171.140 41.590 ;
        RECT 171.360 41.400 172.310 41.680 ;
        RECT 172.480 41.230 172.670 41.670 ;
        RECT 172.840 41.610 173.010 41.840 ;
        RECT 173.180 41.780 173.420 42.180 ;
        RECT 173.590 42.140 174.505 42.440 ;
        RECT 173.590 41.965 173.915 42.140 ;
        RECT 173.590 41.610 173.910 41.965 ;
        RECT 174.675 41.940 174.885 42.590 ;
        RECT 175.525 42.120 175.875 42.770 ;
        RECT 172.840 41.440 173.910 41.610 ;
        RECT 174.155 41.230 174.460 41.690 ;
        RECT 174.630 41.410 174.885 41.940 ;
        RECT 175.060 41.230 175.350 41.955 ;
        RECT 176.045 41.950 176.275 42.940 ;
        RECT 175.525 41.780 176.275 41.950 ;
        RECT 175.525 41.490 175.780 41.780 ;
        RECT 175.950 41.230 176.280 41.610 ;
        RECT 176.450 41.490 176.620 43.610 ;
        RECT 176.790 42.810 177.115 43.595 ;
        RECT 177.285 43.320 177.535 43.780 ;
        RECT 177.705 43.280 177.955 43.610 ;
        RECT 178.170 43.280 178.850 43.610 ;
        RECT 177.705 43.150 177.875 43.280 ;
        RECT 177.480 42.980 177.875 43.150 ;
        RECT 176.850 41.760 177.310 42.810 ;
        RECT 177.480 41.620 177.650 42.980 ;
        RECT 178.045 42.720 178.510 43.110 ;
        RECT 177.820 41.910 178.170 42.530 ;
        RECT 178.340 42.130 178.510 42.720 ;
        RECT 178.680 42.500 178.850 43.280 ;
        RECT 179.020 43.180 179.190 43.520 ;
        RECT 179.425 43.350 179.755 43.780 ;
        RECT 179.925 43.180 180.095 43.520 ;
        RECT 180.390 43.320 180.760 43.780 ;
        RECT 179.020 43.010 180.095 43.180 ;
        RECT 180.930 43.150 181.100 43.610 ;
        RECT 181.335 43.270 182.205 43.610 ;
        RECT 182.375 43.320 182.625 43.780 ;
        RECT 180.540 42.980 181.100 43.150 ;
        RECT 180.540 42.840 180.710 42.980 ;
        RECT 179.210 42.670 180.710 42.840 ;
        RECT 181.405 42.810 181.865 43.100 ;
        RECT 178.680 42.330 180.370 42.500 ;
        RECT 178.340 41.910 178.695 42.130 ;
        RECT 178.865 41.620 179.035 42.330 ;
        RECT 179.240 41.910 180.030 42.160 ;
        RECT 180.200 42.150 180.370 42.330 ;
        RECT 180.540 41.980 180.710 42.670 ;
        RECT 176.980 41.230 177.310 41.590 ;
        RECT 177.480 41.450 177.975 41.620 ;
        RECT 178.180 41.450 179.035 41.620 ;
        RECT 179.910 41.230 180.240 41.690 ;
        RECT 180.450 41.590 180.710 41.980 ;
        RECT 180.900 42.800 181.865 42.810 ;
        RECT 182.035 42.890 182.205 43.270 ;
        RECT 182.795 43.230 182.965 43.520 ;
        RECT 183.145 43.400 183.475 43.780 ;
        RECT 182.795 43.060 183.595 43.230 ;
        RECT 180.900 42.640 181.575 42.800 ;
        RECT 182.035 42.720 183.255 42.890 ;
        RECT 180.900 41.850 181.110 42.640 ;
        RECT 182.035 42.630 182.205 42.720 ;
        RECT 181.280 41.850 181.630 42.470 ;
        RECT 181.800 42.460 182.205 42.630 ;
        RECT 181.800 41.680 181.970 42.460 ;
        RECT 182.140 42.010 182.360 42.290 ;
        RECT 182.540 42.180 183.080 42.550 ;
        RECT 183.425 42.470 183.595 43.060 ;
        RECT 183.815 42.640 184.120 43.780 ;
        RECT 184.290 42.590 184.545 43.470 ;
        RECT 184.720 42.690 186.390 43.780 ;
        RECT 183.425 42.440 184.165 42.470 ;
        RECT 182.140 41.840 182.670 42.010 ;
        RECT 180.450 41.420 180.800 41.590 ;
        RECT 181.020 41.400 181.970 41.680 ;
        RECT 182.140 41.230 182.330 41.670 ;
        RECT 182.500 41.610 182.670 41.840 ;
        RECT 182.840 41.780 183.080 42.180 ;
        RECT 183.250 42.140 184.165 42.440 ;
        RECT 183.250 41.965 183.575 42.140 ;
        RECT 183.250 41.610 183.570 41.965 ;
        RECT 184.335 41.940 184.545 42.590 ;
        RECT 182.500 41.440 183.570 41.610 ;
        RECT 183.815 41.230 184.120 41.690 ;
        RECT 184.290 41.410 184.545 41.940 ;
        RECT 184.720 42.000 185.470 42.520 ;
        RECT 185.640 42.170 186.390 42.690 ;
        RECT 186.610 42.640 186.860 43.780 ;
        RECT 187.030 42.590 187.280 43.470 ;
        RECT 187.450 42.640 187.755 43.780 ;
        RECT 188.095 43.400 188.425 43.780 ;
        RECT 188.605 43.230 188.775 43.520 ;
        RECT 188.945 43.320 189.195 43.780 ;
        RECT 187.975 43.060 188.775 43.230 ;
        RECT 189.365 43.270 190.235 43.610 ;
        RECT 184.720 41.230 186.390 42.000 ;
        RECT 186.610 41.230 186.860 41.985 ;
        RECT 187.030 41.940 187.235 42.590 ;
        RECT 187.975 42.470 188.145 43.060 ;
        RECT 189.365 42.890 189.535 43.270 ;
        RECT 190.470 43.150 190.640 43.610 ;
        RECT 190.810 43.320 191.180 43.780 ;
        RECT 191.475 43.180 191.645 43.520 ;
        RECT 191.815 43.350 192.145 43.780 ;
        RECT 192.380 43.180 192.550 43.520 ;
        RECT 188.315 42.720 189.535 42.890 ;
        RECT 189.705 42.810 190.165 43.100 ;
        RECT 190.470 42.980 191.030 43.150 ;
        RECT 191.475 43.010 192.550 43.180 ;
        RECT 192.720 43.280 193.400 43.610 ;
        RECT 193.615 43.280 193.865 43.610 ;
        RECT 194.035 43.320 194.285 43.780 ;
        RECT 190.860 42.840 191.030 42.980 ;
        RECT 189.705 42.800 190.670 42.810 ;
        RECT 189.365 42.630 189.535 42.720 ;
        RECT 189.995 42.640 190.670 42.800 ;
        RECT 187.405 42.440 188.145 42.470 ;
        RECT 187.405 42.140 188.320 42.440 ;
        RECT 187.995 41.965 188.320 42.140 ;
        RECT 187.030 41.410 187.280 41.940 ;
        RECT 187.450 41.230 187.755 41.690 ;
        RECT 188.000 41.610 188.320 41.965 ;
        RECT 188.490 42.180 189.030 42.550 ;
        RECT 189.365 42.460 189.770 42.630 ;
        RECT 188.490 41.780 188.730 42.180 ;
        RECT 189.210 42.010 189.430 42.290 ;
        RECT 188.900 41.840 189.430 42.010 ;
        RECT 188.900 41.610 189.070 41.840 ;
        RECT 189.600 41.680 189.770 42.460 ;
        RECT 189.940 41.850 190.290 42.470 ;
        RECT 190.460 41.850 190.670 42.640 ;
        RECT 190.860 42.670 192.360 42.840 ;
        RECT 190.860 41.980 191.030 42.670 ;
        RECT 192.720 42.500 192.890 43.280 ;
        RECT 193.695 43.150 193.865 43.280 ;
        RECT 191.200 42.330 192.890 42.500 ;
        RECT 193.060 42.720 193.525 43.110 ;
        RECT 193.695 42.980 194.090 43.150 ;
        RECT 191.200 42.150 191.370 42.330 ;
        RECT 188.000 41.440 189.070 41.610 ;
        RECT 189.240 41.230 189.430 41.670 ;
        RECT 189.600 41.400 190.550 41.680 ;
        RECT 190.860 41.590 191.120 41.980 ;
        RECT 191.540 41.910 192.330 42.160 ;
        RECT 190.770 41.420 191.120 41.590 ;
        RECT 191.330 41.230 191.660 41.690 ;
        RECT 192.535 41.620 192.705 42.330 ;
        RECT 193.060 42.130 193.230 42.720 ;
        RECT 192.875 41.910 193.230 42.130 ;
        RECT 193.400 41.910 193.750 42.530 ;
        RECT 193.920 41.620 194.090 42.980 ;
        RECT 194.455 42.810 194.780 43.595 ;
        RECT 194.260 41.760 194.720 42.810 ;
        RECT 192.535 41.450 193.390 41.620 ;
        RECT 193.595 41.450 194.090 41.620 ;
        RECT 194.260 41.230 194.590 41.590 ;
        RECT 194.950 41.490 195.120 43.610 ;
        RECT 195.290 43.280 195.620 43.780 ;
        RECT 195.790 43.110 196.045 43.610 ;
        RECT 195.295 42.940 196.045 43.110 ;
        RECT 195.295 41.950 195.525 42.940 ;
        RECT 195.695 42.120 196.045 42.770 ;
        RECT 196.220 42.690 199.730 43.780 ;
        RECT 196.220 42.000 197.870 42.520 ;
        RECT 198.040 42.170 199.730 42.690 ;
        RECT 200.820 42.615 201.110 43.780 ;
        RECT 201.285 43.110 201.540 43.610 ;
        RECT 201.710 43.280 202.040 43.780 ;
        RECT 201.285 42.940 202.035 43.110 ;
        RECT 201.285 42.120 201.635 42.770 ;
        RECT 195.295 41.780 196.045 41.950 ;
        RECT 195.290 41.230 195.620 41.610 ;
        RECT 195.790 41.490 196.045 41.780 ;
        RECT 196.220 41.230 199.730 42.000 ;
        RECT 200.820 41.230 201.110 41.955 ;
        RECT 201.805 41.950 202.035 42.940 ;
        RECT 201.285 41.780 202.035 41.950 ;
        RECT 201.285 41.490 201.540 41.780 ;
        RECT 201.710 41.230 202.040 41.610 ;
        RECT 202.210 41.490 202.380 43.610 ;
        RECT 202.550 42.810 202.875 43.595 ;
        RECT 203.045 43.320 203.295 43.780 ;
        RECT 203.465 43.280 203.715 43.610 ;
        RECT 203.930 43.280 204.610 43.610 ;
        RECT 203.465 43.150 203.635 43.280 ;
        RECT 203.240 42.980 203.635 43.150 ;
        RECT 202.610 41.760 203.070 42.810 ;
        RECT 203.240 41.620 203.410 42.980 ;
        RECT 203.805 42.720 204.270 43.110 ;
        RECT 203.580 41.910 203.930 42.530 ;
        RECT 204.100 42.130 204.270 42.720 ;
        RECT 204.440 42.500 204.610 43.280 ;
        RECT 204.780 43.180 204.950 43.520 ;
        RECT 205.185 43.350 205.515 43.780 ;
        RECT 205.685 43.180 205.855 43.520 ;
        RECT 206.150 43.320 206.520 43.780 ;
        RECT 204.780 43.010 205.855 43.180 ;
        RECT 206.690 43.150 206.860 43.610 ;
        RECT 207.095 43.270 207.965 43.610 ;
        RECT 208.135 43.320 208.385 43.780 ;
        RECT 206.300 42.980 206.860 43.150 ;
        RECT 206.300 42.840 206.470 42.980 ;
        RECT 204.970 42.670 206.470 42.840 ;
        RECT 207.165 42.810 207.625 43.100 ;
        RECT 204.440 42.330 206.130 42.500 ;
        RECT 204.100 41.910 204.455 42.130 ;
        RECT 204.625 41.620 204.795 42.330 ;
        RECT 205.000 41.910 205.790 42.160 ;
        RECT 205.960 42.150 206.130 42.330 ;
        RECT 206.300 41.980 206.470 42.670 ;
        RECT 202.740 41.230 203.070 41.590 ;
        RECT 203.240 41.450 203.735 41.620 ;
        RECT 203.940 41.450 204.795 41.620 ;
        RECT 205.670 41.230 206.000 41.690 ;
        RECT 206.210 41.590 206.470 41.980 ;
        RECT 206.660 42.800 207.625 42.810 ;
        RECT 207.795 42.890 207.965 43.270 ;
        RECT 208.555 43.230 208.725 43.520 ;
        RECT 208.905 43.400 209.235 43.780 ;
        RECT 208.555 43.060 209.355 43.230 ;
        RECT 206.660 42.640 207.335 42.800 ;
        RECT 207.795 42.720 209.015 42.890 ;
        RECT 206.660 41.850 206.870 42.640 ;
        RECT 207.795 42.630 207.965 42.720 ;
        RECT 207.040 41.850 207.390 42.470 ;
        RECT 207.560 42.460 207.965 42.630 ;
        RECT 207.560 41.680 207.730 42.460 ;
        RECT 207.900 42.010 208.120 42.290 ;
        RECT 208.300 42.180 208.840 42.550 ;
        RECT 209.185 42.470 209.355 43.060 ;
        RECT 209.575 42.640 209.880 43.780 ;
        RECT 210.050 42.590 210.305 43.470 ;
        RECT 209.185 42.440 209.925 42.470 ;
        RECT 207.900 41.840 208.430 42.010 ;
        RECT 206.210 41.420 206.560 41.590 ;
        RECT 206.780 41.400 207.730 41.680 ;
        RECT 207.900 41.230 208.090 41.670 ;
        RECT 208.260 41.610 208.430 41.840 ;
        RECT 208.600 41.780 208.840 42.180 ;
        RECT 209.010 42.140 209.925 42.440 ;
        RECT 209.010 41.965 209.335 42.140 ;
        RECT 209.010 41.610 209.330 41.965 ;
        RECT 210.095 41.940 210.305 42.590 ;
        RECT 208.260 41.440 209.330 41.610 ;
        RECT 209.575 41.230 209.880 41.690 ;
        RECT 210.050 41.410 210.305 41.940 ;
        RECT 210.480 42.640 210.865 43.610 ;
        RECT 211.035 43.320 211.360 43.780 ;
        RECT 211.880 43.150 212.160 43.610 ;
        RECT 211.035 42.930 212.160 43.150 ;
        RECT 210.480 41.970 210.760 42.640 ;
        RECT 211.035 42.470 211.485 42.930 ;
        RECT 212.350 42.760 212.750 43.610 ;
        RECT 213.150 43.320 213.420 43.780 ;
        RECT 213.590 43.150 213.875 43.610 ;
        RECT 210.930 42.140 211.485 42.470 ;
        RECT 211.655 42.200 212.750 42.760 ;
        RECT 211.035 42.030 211.485 42.140 ;
        RECT 210.480 41.400 210.865 41.970 ;
        RECT 211.035 41.860 212.160 42.030 ;
        RECT 211.035 41.230 211.360 41.690 ;
        RECT 211.880 41.400 212.160 41.860 ;
        RECT 212.350 41.400 212.750 42.200 ;
        RECT 212.920 42.930 213.875 43.150 ;
        RECT 215.085 43.110 215.340 43.610 ;
        RECT 215.510 43.280 215.840 43.780 ;
        RECT 215.085 42.940 215.835 43.110 ;
        RECT 212.920 42.030 213.130 42.930 ;
        RECT 213.300 42.200 213.990 42.760 ;
        RECT 215.085 42.120 215.435 42.770 ;
        RECT 212.920 41.860 213.875 42.030 ;
        RECT 215.605 41.950 215.835 42.940 ;
        RECT 213.150 41.230 213.420 41.690 ;
        RECT 213.590 41.400 213.875 41.860 ;
        RECT 215.085 41.780 215.835 41.950 ;
        RECT 215.085 41.490 215.340 41.780 ;
        RECT 215.510 41.230 215.840 41.610 ;
        RECT 216.010 41.490 216.180 43.610 ;
        RECT 216.350 42.810 216.675 43.595 ;
        RECT 216.845 43.320 217.095 43.780 ;
        RECT 217.265 43.280 217.515 43.610 ;
        RECT 217.730 43.280 218.410 43.610 ;
        RECT 217.265 43.150 217.435 43.280 ;
        RECT 217.040 42.980 217.435 43.150 ;
        RECT 216.410 41.760 216.870 42.810 ;
        RECT 217.040 41.620 217.210 42.980 ;
        RECT 217.605 42.720 218.070 43.110 ;
        RECT 217.380 41.910 217.730 42.530 ;
        RECT 217.900 42.130 218.070 42.720 ;
        RECT 218.240 42.500 218.410 43.280 ;
        RECT 218.580 43.180 218.750 43.520 ;
        RECT 218.985 43.350 219.315 43.780 ;
        RECT 219.485 43.180 219.655 43.520 ;
        RECT 219.950 43.320 220.320 43.780 ;
        RECT 218.580 43.010 219.655 43.180 ;
        RECT 220.490 43.150 220.660 43.610 ;
        RECT 220.895 43.270 221.765 43.610 ;
        RECT 221.935 43.320 222.185 43.780 ;
        RECT 220.100 42.980 220.660 43.150 ;
        RECT 220.100 42.840 220.270 42.980 ;
        RECT 218.770 42.670 220.270 42.840 ;
        RECT 220.965 42.810 221.425 43.100 ;
        RECT 218.240 42.330 219.930 42.500 ;
        RECT 217.900 41.910 218.255 42.130 ;
        RECT 218.425 41.620 218.595 42.330 ;
        RECT 218.800 41.910 219.590 42.160 ;
        RECT 219.760 42.150 219.930 42.330 ;
        RECT 220.100 41.980 220.270 42.670 ;
        RECT 216.540 41.230 216.870 41.590 ;
        RECT 217.040 41.450 217.535 41.620 ;
        RECT 217.740 41.450 218.595 41.620 ;
        RECT 219.470 41.230 219.800 41.690 ;
        RECT 220.010 41.590 220.270 41.980 ;
        RECT 220.460 42.800 221.425 42.810 ;
        RECT 221.595 42.890 221.765 43.270 ;
        RECT 222.355 43.230 222.525 43.520 ;
        RECT 222.705 43.400 223.035 43.780 ;
        RECT 222.355 43.060 223.155 43.230 ;
        RECT 220.460 42.640 221.135 42.800 ;
        RECT 221.595 42.720 222.815 42.890 ;
        RECT 220.460 41.850 220.670 42.640 ;
        RECT 221.595 42.630 221.765 42.720 ;
        RECT 220.840 41.850 221.190 42.470 ;
        RECT 221.360 42.460 221.765 42.630 ;
        RECT 221.360 41.680 221.530 42.460 ;
        RECT 221.700 42.010 221.920 42.290 ;
        RECT 222.100 42.180 222.640 42.550 ;
        RECT 222.985 42.470 223.155 43.060 ;
        RECT 223.375 42.640 223.680 43.780 ;
        RECT 223.850 42.590 224.100 43.470 ;
        RECT 224.270 42.640 224.520 43.780 ;
        RECT 224.740 42.690 226.410 43.780 ;
        RECT 222.985 42.440 223.725 42.470 ;
        RECT 221.700 41.840 222.230 42.010 ;
        RECT 220.010 41.420 220.360 41.590 ;
        RECT 220.580 41.400 221.530 41.680 ;
        RECT 221.700 41.230 221.890 41.670 ;
        RECT 222.060 41.610 222.230 41.840 ;
        RECT 222.400 41.780 222.640 42.180 ;
        RECT 222.810 42.140 223.725 42.440 ;
        RECT 222.810 41.965 223.135 42.140 ;
        RECT 222.810 41.610 223.130 41.965 ;
        RECT 223.895 41.940 224.100 42.590 ;
        RECT 224.740 42.000 225.490 42.520 ;
        RECT 225.660 42.170 226.410 42.690 ;
        RECT 226.580 42.615 226.870 43.780 ;
        RECT 227.095 42.910 227.380 43.780 ;
        RECT 227.550 43.150 227.810 43.610 ;
        RECT 227.985 43.320 228.240 43.780 ;
        RECT 228.410 43.150 228.670 43.610 ;
        RECT 227.550 42.980 228.670 43.150 ;
        RECT 228.840 42.980 229.150 43.780 ;
        RECT 227.550 42.730 227.810 42.980 ;
        RECT 229.320 42.810 229.630 43.610 ;
        RECT 227.055 42.560 227.810 42.730 ;
        RECT 228.600 42.640 229.630 42.810 ;
        RECT 227.055 42.050 227.460 42.560 ;
        RECT 228.600 42.390 228.770 42.640 ;
        RECT 227.630 42.220 228.770 42.390 ;
        RECT 222.060 41.440 223.130 41.610 ;
        RECT 223.375 41.230 223.680 41.690 ;
        RECT 223.850 41.410 224.100 41.940 ;
        RECT 224.270 41.230 224.520 41.985 ;
        RECT 224.740 41.230 226.410 42.000 ;
        RECT 226.580 41.230 226.870 41.955 ;
        RECT 227.055 41.880 228.705 42.050 ;
        RECT 228.940 41.900 229.290 42.470 ;
        RECT 227.100 41.230 227.380 41.710 ;
        RECT 227.550 41.490 227.810 41.880 ;
        RECT 227.985 41.230 228.240 41.710 ;
        RECT 228.410 41.490 228.705 41.880 ;
        RECT 229.460 41.730 229.630 42.640 ;
        RECT 228.885 41.230 229.160 41.710 ;
        RECT 229.330 41.400 229.630 41.730 ;
        RECT 230.720 42.640 231.105 43.610 ;
        RECT 231.275 43.320 231.600 43.780 ;
        RECT 232.120 43.150 232.400 43.610 ;
        RECT 231.275 42.930 232.400 43.150 ;
        RECT 230.720 41.970 231.000 42.640 ;
        RECT 231.275 42.470 231.725 42.930 ;
        RECT 232.590 42.760 232.990 43.610 ;
        RECT 233.390 43.320 233.660 43.780 ;
        RECT 233.830 43.150 234.115 43.610 ;
        RECT 231.170 42.140 231.725 42.470 ;
        RECT 231.895 42.200 232.990 42.760 ;
        RECT 231.275 42.030 231.725 42.140 ;
        RECT 230.720 41.400 231.105 41.970 ;
        RECT 231.275 41.860 232.400 42.030 ;
        RECT 231.275 41.230 231.600 41.690 ;
        RECT 232.120 41.400 232.400 41.860 ;
        RECT 232.590 41.400 232.990 42.200 ;
        RECT 233.160 42.930 234.115 43.150 ;
        RECT 234.860 43.020 235.525 43.610 ;
        RECT 233.160 42.030 233.370 42.930 ;
        RECT 233.540 42.200 234.230 42.760 ;
        RECT 234.860 42.050 235.110 43.020 ;
        RECT 235.695 42.940 236.025 43.780 ;
        RECT 236.535 43.190 237.340 43.610 ;
        RECT 236.195 43.020 237.760 43.190 ;
        RECT 236.195 42.770 236.365 43.020 ;
        RECT 235.445 42.600 236.365 42.770 ;
        RECT 236.535 42.760 236.910 42.850 ;
        RECT 235.445 42.430 235.615 42.600 ;
        RECT 236.535 42.590 236.930 42.760 ;
        RECT 236.535 42.430 236.910 42.590 ;
        RECT 235.280 42.220 235.615 42.430 ;
        RECT 235.785 42.220 236.235 42.430 ;
        RECT 236.425 42.220 236.910 42.430 ;
        RECT 237.100 42.470 237.420 42.850 ;
        RECT 237.590 42.770 237.760 43.020 ;
        RECT 237.930 42.940 238.180 43.780 ;
        RECT 238.375 42.770 238.675 43.610 ;
        RECT 237.590 42.600 238.675 42.770 ;
        RECT 239.000 42.690 240.210 43.780 ;
        RECT 237.100 42.220 237.480 42.470 ;
        RECT 237.660 42.220 237.990 42.430 ;
        RECT 233.160 41.860 234.115 42.030 ;
        RECT 233.390 41.230 233.660 41.690 ;
        RECT 233.830 41.400 234.115 41.860 ;
        RECT 234.860 41.410 235.545 42.050 ;
        RECT 235.715 41.230 235.885 42.050 ;
        RECT 236.055 41.880 237.755 42.050 ;
        RECT 236.055 41.415 236.385 41.880 ;
        RECT 237.370 41.790 237.755 41.880 ;
        RECT 238.160 41.970 238.330 42.600 ;
        RECT 238.500 42.140 238.830 42.430 ;
        RECT 239.000 41.980 239.520 42.520 ;
        RECT 239.690 42.150 240.210 42.690 ;
        RECT 240.385 42.640 240.720 43.610 ;
        RECT 240.890 42.640 241.060 43.780 ;
        RECT 241.230 43.440 243.260 43.610 ;
        RECT 238.160 41.790 238.670 41.970 ;
        RECT 236.555 41.230 236.725 41.700 ;
        RECT 236.985 41.450 238.170 41.620 ;
        RECT 238.340 41.400 238.670 41.790 ;
        RECT 239.000 41.230 240.210 41.980 ;
        RECT 240.385 41.970 240.555 42.640 ;
        RECT 241.230 42.470 241.400 43.440 ;
        RECT 240.725 42.140 240.980 42.470 ;
        RECT 241.205 42.140 241.400 42.470 ;
        RECT 241.570 43.100 242.695 43.270 ;
        RECT 240.810 41.970 240.980 42.140 ;
        RECT 241.570 41.970 241.740 43.100 ;
        RECT 240.385 41.400 240.640 41.970 ;
        RECT 240.810 41.800 241.740 41.970 ;
        RECT 241.910 42.760 242.920 42.930 ;
        RECT 241.910 41.960 242.080 42.760 ;
        RECT 241.565 41.765 241.740 41.800 ;
        RECT 240.810 41.230 241.140 41.630 ;
        RECT 241.565 41.400 242.095 41.765 ;
        RECT 242.285 41.740 242.560 42.560 ;
        RECT 242.280 41.570 242.560 41.740 ;
        RECT 242.285 41.400 242.560 41.570 ;
        RECT 242.730 41.400 242.920 42.760 ;
        RECT 243.090 42.775 243.260 43.440 ;
        RECT 243.430 43.020 243.600 43.780 ;
        RECT 243.835 43.020 244.350 43.430 ;
        RECT 243.090 42.585 243.840 42.775 ;
        RECT 244.010 42.210 244.350 43.020 ;
        RECT 244.635 43.150 244.920 43.610 ;
        RECT 245.090 43.320 245.360 43.780 ;
        RECT 244.635 42.930 245.590 43.150 ;
        RECT 243.120 42.040 244.350 42.210 ;
        RECT 244.520 42.200 245.210 42.760 ;
        RECT 243.100 41.230 243.610 41.765 ;
        RECT 243.830 41.435 244.075 42.040 ;
        RECT 245.380 42.030 245.590 42.930 ;
        RECT 244.635 41.860 245.590 42.030 ;
        RECT 245.760 42.760 246.160 43.610 ;
        RECT 246.350 43.150 246.630 43.610 ;
        RECT 247.150 43.320 247.475 43.780 ;
        RECT 246.350 42.930 247.475 43.150 ;
        RECT 245.760 42.200 246.855 42.760 ;
        RECT 247.025 42.470 247.475 42.930 ;
        RECT 247.645 42.640 248.030 43.610 ;
        RECT 244.635 41.400 244.920 41.860 ;
        RECT 245.090 41.230 245.360 41.690 ;
        RECT 245.760 41.400 246.160 42.200 ;
        RECT 247.025 42.140 247.580 42.470 ;
        RECT 247.025 42.030 247.475 42.140 ;
        RECT 246.350 41.860 247.475 42.030 ;
        RECT 247.750 41.970 248.030 42.640 ;
        RECT 246.350 41.400 246.630 41.860 ;
        RECT 247.150 41.230 247.475 41.690 ;
        RECT 247.645 41.400 248.030 41.970 ;
        RECT 248.235 42.990 248.770 43.610 ;
        RECT 248.235 41.970 248.550 42.990 ;
        RECT 248.940 42.980 249.270 43.780 ;
        RECT 249.755 42.810 250.145 42.985 ;
        RECT 248.720 42.640 250.145 42.810 ;
        RECT 250.500 42.690 252.170 43.780 ;
        RECT 248.720 42.140 248.890 42.640 ;
        RECT 248.235 41.400 248.850 41.970 ;
        RECT 249.140 41.910 249.405 42.470 ;
        RECT 249.575 41.740 249.745 42.640 ;
        RECT 249.915 41.910 250.270 42.470 ;
        RECT 250.500 42.000 251.250 42.520 ;
        RECT 251.420 42.170 252.170 42.690 ;
        RECT 252.340 42.615 252.630 43.780 ;
        RECT 252.800 42.945 253.145 43.780 ;
        RECT 253.320 42.775 253.575 43.580 ;
        RECT 253.745 42.945 254.005 43.780 ;
        RECT 254.180 42.775 254.435 43.580 ;
        RECT 254.605 42.945 254.865 43.780 ;
        RECT 255.035 42.775 255.295 43.580 ;
        RECT 255.465 42.945 255.850 43.780 ;
        RECT 256.055 42.990 256.590 43.610 ;
        RECT 252.820 42.605 255.850 42.775 ;
        RECT 252.820 42.040 252.990 42.605 ;
        RECT 253.160 42.210 255.375 42.435 ;
        RECT 255.550 42.040 255.850 42.605 ;
        RECT 249.020 41.230 249.235 41.740 ;
        RECT 249.465 41.410 249.745 41.740 ;
        RECT 249.925 41.230 250.165 41.740 ;
        RECT 250.500 41.230 252.170 42.000 ;
        RECT 252.340 41.230 252.630 41.955 ;
        RECT 252.820 41.870 255.850 42.040 ;
        RECT 256.055 41.970 256.370 42.990 ;
        RECT 256.760 42.980 257.090 43.780 ;
        RECT 257.575 42.810 257.965 42.985 ;
        RECT 256.540 42.640 257.965 42.810 ;
        RECT 259.240 42.640 259.520 43.780 ;
        RECT 256.540 42.140 256.710 42.640 ;
        RECT 253.280 41.230 253.575 41.700 ;
        RECT 253.745 41.425 254.005 41.870 ;
        RECT 254.175 41.230 254.435 41.700 ;
        RECT 254.605 41.425 254.860 41.870 ;
        RECT 255.030 41.230 255.330 41.700 ;
        RECT 256.055 41.400 256.670 41.970 ;
        RECT 256.960 41.910 257.225 42.470 ;
        RECT 257.395 41.740 257.565 42.640 ;
        RECT 259.690 42.630 260.020 43.610 ;
        RECT 260.190 42.640 260.450 43.780 ;
        RECT 260.620 42.690 264.130 43.780 ;
        RECT 264.300 42.690 265.510 43.780 ;
        RECT 265.685 43.110 265.940 43.610 ;
        RECT 266.110 43.280 266.440 43.780 ;
        RECT 265.685 42.940 266.435 43.110 ;
        RECT 257.735 41.910 258.090 42.470 ;
        RECT 259.250 42.200 259.585 42.470 ;
        RECT 259.755 42.030 259.925 42.630 ;
        RECT 260.095 42.220 260.430 42.470 ;
        RECT 256.840 41.230 257.055 41.740 ;
        RECT 257.285 41.410 257.565 41.740 ;
        RECT 257.745 41.230 257.985 41.740 ;
        RECT 259.240 41.230 259.550 42.030 ;
        RECT 259.755 41.400 260.450 42.030 ;
        RECT 260.620 42.000 262.270 42.520 ;
        RECT 262.440 42.170 264.130 42.690 ;
        RECT 260.620 41.230 264.130 42.000 ;
        RECT 264.300 41.980 264.820 42.520 ;
        RECT 264.990 42.150 265.510 42.690 ;
        RECT 265.685 42.120 266.035 42.770 ;
        RECT 264.300 41.230 265.510 41.980 ;
        RECT 266.205 41.950 266.435 42.940 ;
        RECT 265.685 41.780 266.435 41.950 ;
        RECT 265.685 41.490 265.940 41.780 ;
        RECT 266.110 41.230 266.440 41.610 ;
        RECT 266.610 41.490 266.780 43.610 ;
        RECT 266.950 42.810 267.275 43.595 ;
        RECT 267.445 43.320 267.695 43.780 ;
        RECT 267.865 43.280 268.115 43.610 ;
        RECT 268.330 43.280 269.010 43.610 ;
        RECT 267.865 43.150 268.035 43.280 ;
        RECT 267.640 42.980 268.035 43.150 ;
        RECT 267.010 41.760 267.470 42.810 ;
        RECT 267.640 41.620 267.810 42.980 ;
        RECT 268.205 42.720 268.670 43.110 ;
        RECT 267.980 41.910 268.330 42.530 ;
        RECT 268.500 42.130 268.670 42.720 ;
        RECT 268.840 42.500 269.010 43.280 ;
        RECT 269.180 43.180 269.350 43.520 ;
        RECT 269.585 43.350 269.915 43.780 ;
        RECT 270.085 43.180 270.255 43.520 ;
        RECT 270.550 43.320 270.920 43.780 ;
        RECT 269.180 43.010 270.255 43.180 ;
        RECT 271.090 43.150 271.260 43.610 ;
        RECT 271.495 43.270 272.365 43.610 ;
        RECT 272.535 43.320 272.785 43.780 ;
        RECT 270.700 42.980 271.260 43.150 ;
        RECT 270.700 42.840 270.870 42.980 ;
        RECT 269.370 42.670 270.870 42.840 ;
        RECT 271.565 42.810 272.025 43.100 ;
        RECT 268.840 42.330 270.530 42.500 ;
        RECT 268.500 41.910 268.855 42.130 ;
        RECT 269.025 41.620 269.195 42.330 ;
        RECT 269.400 41.910 270.190 42.160 ;
        RECT 270.360 42.150 270.530 42.330 ;
        RECT 270.700 41.980 270.870 42.670 ;
        RECT 267.140 41.230 267.470 41.590 ;
        RECT 267.640 41.450 268.135 41.620 ;
        RECT 268.340 41.450 269.195 41.620 ;
        RECT 270.070 41.230 270.400 41.690 ;
        RECT 270.610 41.590 270.870 41.980 ;
        RECT 271.060 42.800 272.025 42.810 ;
        RECT 272.195 42.890 272.365 43.270 ;
        RECT 272.955 43.230 273.125 43.520 ;
        RECT 273.305 43.400 273.635 43.780 ;
        RECT 272.955 43.060 273.755 43.230 ;
        RECT 271.060 42.640 271.735 42.800 ;
        RECT 272.195 42.720 273.415 42.890 ;
        RECT 271.060 41.850 271.270 42.640 ;
        RECT 272.195 42.630 272.365 42.720 ;
        RECT 271.440 41.850 271.790 42.470 ;
        RECT 271.960 42.460 272.365 42.630 ;
        RECT 271.960 41.680 272.130 42.460 ;
        RECT 272.300 42.010 272.520 42.290 ;
        RECT 272.700 42.180 273.240 42.550 ;
        RECT 273.585 42.470 273.755 43.060 ;
        RECT 273.975 42.640 274.280 43.780 ;
        RECT 274.450 42.590 274.705 43.470 ;
        RECT 274.935 42.910 275.220 43.780 ;
        RECT 275.390 43.150 275.650 43.610 ;
        RECT 275.825 43.320 276.080 43.780 ;
        RECT 276.250 43.150 276.510 43.610 ;
        RECT 275.390 42.980 276.510 43.150 ;
        RECT 276.680 42.980 276.990 43.780 ;
        RECT 275.390 42.730 275.650 42.980 ;
        RECT 277.160 42.810 277.470 43.610 ;
        RECT 273.585 42.440 274.325 42.470 ;
        RECT 272.300 41.840 272.830 42.010 ;
        RECT 270.610 41.420 270.960 41.590 ;
        RECT 271.180 41.400 272.130 41.680 ;
        RECT 272.300 41.230 272.490 41.670 ;
        RECT 272.660 41.610 272.830 41.840 ;
        RECT 273.000 41.780 273.240 42.180 ;
        RECT 273.410 42.140 274.325 42.440 ;
        RECT 273.410 41.965 273.735 42.140 ;
        RECT 273.410 41.610 273.730 41.965 ;
        RECT 274.495 41.940 274.705 42.590 ;
        RECT 272.660 41.440 273.730 41.610 ;
        RECT 273.975 41.230 274.280 41.690 ;
        RECT 274.450 41.410 274.705 41.940 ;
        RECT 274.895 42.560 275.650 42.730 ;
        RECT 276.440 42.640 277.470 42.810 ;
        RECT 274.895 42.050 275.300 42.560 ;
        RECT 276.440 42.390 276.610 42.640 ;
        RECT 275.470 42.220 276.610 42.390 ;
        RECT 274.895 41.880 276.545 42.050 ;
        RECT 276.780 41.900 277.130 42.470 ;
        RECT 274.940 41.230 275.220 41.710 ;
        RECT 275.390 41.490 275.650 41.880 ;
        RECT 275.825 41.230 276.080 41.710 ;
        RECT 276.250 41.490 276.545 41.880 ;
        RECT 277.300 41.730 277.470 42.640 ;
        RECT 278.100 42.615 278.390 43.780 ;
        RECT 278.560 42.640 278.945 43.610 ;
        RECT 279.115 43.320 279.440 43.780 ;
        RECT 279.960 43.150 280.240 43.610 ;
        RECT 279.115 42.930 280.240 43.150 ;
        RECT 278.560 41.970 278.840 42.640 ;
        RECT 279.115 42.470 279.565 42.930 ;
        RECT 280.430 42.760 280.830 43.610 ;
        RECT 281.230 43.320 281.500 43.780 ;
        RECT 281.670 43.150 281.955 43.610 ;
        RECT 279.010 42.140 279.565 42.470 ;
        RECT 279.735 42.200 280.830 42.760 ;
        RECT 279.115 42.030 279.565 42.140 ;
        RECT 276.725 41.230 277.000 41.710 ;
        RECT 277.170 41.400 277.470 41.730 ;
        RECT 278.100 41.230 278.390 41.955 ;
        RECT 278.560 41.400 278.945 41.970 ;
        RECT 279.115 41.860 280.240 42.030 ;
        RECT 279.115 41.230 279.440 41.690 ;
        RECT 279.960 41.400 280.240 41.860 ;
        RECT 280.430 41.400 280.830 42.200 ;
        RECT 281.000 42.930 281.955 43.150 ;
        RECT 281.000 42.030 281.210 42.930 ;
        RECT 281.380 42.200 282.070 42.760 ;
        RECT 282.240 42.690 284.830 43.780 ;
        RECT 281.000 41.860 281.955 42.030 ;
        RECT 281.230 41.230 281.500 41.690 ;
        RECT 281.670 41.400 281.955 41.860 ;
        RECT 282.240 42.000 283.450 42.520 ;
        RECT 283.620 42.170 284.830 42.690 ;
        RECT 285.465 42.590 285.720 43.470 ;
        RECT 285.890 42.640 286.195 43.780 ;
        RECT 286.535 43.400 286.865 43.780 ;
        RECT 287.045 43.230 287.215 43.520 ;
        RECT 287.385 43.320 287.635 43.780 ;
        RECT 286.415 43.060 287.215 43.230 ;
        RECT 287.805 43.270 288.675 43.610 ;
        RECT 282.240 41.230 284.830 42.000 ;
        RECT 285.465 41.940 285.675 42.590 ;
        RECT 286.415 42.470 286.585 43.060 ;
        RECT 287.805 42.890 287.975 43.270 ;
        RECT 288.910 43.150 289.080 43.610 ;
        RECT 289.250 43.320 289.620 43.780 ;
        RECT 289.915 43.180 290.085 43.520 ;
        RECT 290.255 43.350 290.585 43.780 ;
        RECT 290.820 43.180 290.990 43.520 ;
        RECT 286.755 42.720 287.975 42.890 ;
        RECT 288.145 42.810 288.605 43.100 ;
        RECT 288.910 42.980 289.470 43.150 ;
        RECT 289.915 43.010 290.990 43.180 ;
        RECT 291.160 43.280 291.840 43.610 ;
        RECT 292.055 43.280 292.305 43.610 ;
        RECT 292.475 43.320 292.725 43.780 ;
        RECT 289.300 42.840 289.470 42.980 ;
        RECT 288.145 42.800 289.110 42.810 ;
        RECT 287.805 42.630 287.975 42.720 ;
        RECT 288.435 42.640 289.110 42.800 ;
        RECT 285.845 42.440 286.585 42.470 ;
        RECT 285.845 42.140 286.760 42.440 ;
        RECT 286.435 41.965 286.760 42.140 ;
        RECT 285.465 41.410 285.720 41.940 ;
        RECT 285.890 41.230 286.195 41.690 ;
        RECT 286.440 41.610 286.760 41.965 ;
        RECT 286.930 42.180 287.470 42.550 ;
        RECT 287.805 42.460 288.210 42.630 ;
        RECT 286.930 41.780 287.170 42.180 ;
        RECT 287.650 42.010 287.870 42.290 ;
        RECT 287.340 41.840 287.870 42.010 ;
        RECT 287.340 41.610 287.510 41.840 ;
        RECT 288.040 41.680 288.210 42.460 ;
        RECT 288.380 41.850 288.730 42.470 ;
        RECT 288.900 41.850 289.110 42.640 ;
        RECT 289.300 42.670 290.800 42.840 ;
        RECT 289.300 41.980 289.470 42.670 ;
        RECT 291.160 42.500 291.330 43.280 ;
        RECT 292.135 43.150 292.305 43.280 ;
        RECT 289.640 42.330 291.330 42.500 ;
        RECT 291.500 42.720 291.965 43.110 ;
        RECT 292.135 42.980 292.530 43.150 ;
        RECT 289.640 42.150 289.810 42.330 ;
        RECT 286.440 41.440 287.510 41.610 ;
        RECT 287.680 41.230 287.870 41.670 ;
        RECT 288.040 41.400 288.990 41.680 ;
        RECT 289.300 41.590 289.560 41.980 ;
        RECT 289.980 41.910 290.770 42.160 ;
        RECT 289.210 41.420 289.560 41.590 ;
        RECT 289.770 41.230 290.100 41.690 ;
        RECT 290.975 41.620 291.145 42.330 ;
        RECT 291.500 42.130 291.670 42.720 ;
        RECT 291.315 41.910 291.670 42.130 ;
        RECT 291.840 41.910 292.190 42.530 ;
        RECT 292.360 41.620 292.530 42.980 ;
        RECT 292.895 42.810 293.220 43.595 ;
        RECT 292.700 41.760 293.160 42.810 ;
        RECT 290.975 41.450 291.830 41.620 ;
        RECT 292.035 41.450 292.530 41.620 ;
        RECT 292.700 41.230 293.030 41.590 ;
        RECT 293.390 41.490 293.560 43.610 ;
        RECT 293.730 43.280 294.060 43.780 ;
        RECT 294.230 43.110 294.485 43.610 ;
        RECT 294.660 43.345 300.005 43.780 ;
        RECT 293.735 42.940 294.485 43.110 ;
        RECT 293.735 41.950 293.965 42.940 ;
        RECT 294.135 42.120 294.485 42.770 ;
        RECT 293.735 41.780 294.485 41.950 ;
        RECT 293.730 41.230 294.060 41.610 ;
        RECT 294.230 41.490 294.485 41.780 ;
        RECT 296.245 41.775 296.585 42.605 ;
        RECT 298.065 42.095 298.415 43.345 ;
        RECT 300.180 42.690 303.690 43.780 ;
        RECT 300.180 42.000 301.830 42.520 ;
        RECT 302.000 42.170 303.690 42.690 ;
        RECT 303.860 42.615 304.150 43.780 ;
        RECT 304.320 42.810 304.590 43.580 ;
        RECT 304.760 43.000 305.090 43.780 ;
        RECT 305.295 43.175 305.480 43.580 ;
        RECT 305.650 43.355 305.985 43.780 ;
        RECT 305.295 43.000 305.960 43.175 ;
        RECT 304.320 42.640 305.450 42.810 ;
        RECT 294.660 41.230 300.005 41.775 ;
        RECT 300.180 41.230 303.690 42.000 ;
        RECT 303.860 41.230 304.150 41.955 ;
        RECT 304.320 41.730 304.490 42.640 ;
        RECT 304.660 41.890 305.020 42.470 ;
        RECT 305.200 42.140 305.450 42.640 ;
        RECT 305.620 41.970 305.960 43.000 ;
        RECT 306.275 43.150 306.560 43.610 ;
        RECT 306.730 43.320 307.000 43.780 ;
        RECT 306.275 42.930 307.230 43.150 ;
        RECT 306.160 42.200 306.850 42.760 ;
        RECT 307.020 42.030 307.230 42.930 ;
        RECT 305.275 41.800 305.960 41.970 ;
        RECT 306.275 41.860 307.230 42.030 ;
        RECT 307.400 42.760 307.800 43.610 ;
        RECT 307.990 43.150 308.270 43.610 ;
        RECT 308.790 43.320 309.115 43.780 ;
        RECT 307.990 42.930 309.115 43.150 ;
        RECT 307.400 42.200 308.495 42.760 ;
        RECT 308.665 42.470 309.115 42.930 ;
        RECT 309.285 42.640 309.670 43.610 ;
        RECT 304.320 41.400 304.580 41.730 ;
        RECT 304.790 41.230 305.065 41.710 ;
        RECT 305.275 41.400 305.480 41.800 ;
        RECT 305.650 41.230 305.985 41.630 ;
        RECT 306.275 41.400 306.560 41.860 ;
        RECT 306.730 41.230 307.000 41.690 ;
        RECT 307.400 41.400 307.800 42.200 ;
        RECT 308.665 42.140 309.220 42.470 ;
        RECT 308.665 42.030 309.115 42.140 ;
        RECT 307.990 41.860 309.115 42.030 ;
        RECT 309.390 41.970 309.670 42.640 ;
        RECT 309.840 42.690 311.050 43.780 ;
        RECT 309.840 42.150 310.360 42.690 ;
        RECT 310.530 41.980 311.050 42.520 ;
        RECT 307.990 41.400 308.270 41.860 ;
        RECT 308.790 41.230 309.115 41.690 ;
        RECT 309.285 41.400 309.670 41.970 ;
        RECT 309.840 41.230 311.050 41.980 ;
        RECT 162.095 41.060 311.135 41.230 ;
        RECT 162.180 40.310 163.390 41.060 ;
        RECT 162.180 39.770 162.700 40.310 ;
        RECT 163.560 40.290 167.070 41.060 ;
        RECT 168.165 40.510 168.420 40.800 ;
        RECT 168.590 40.680 168.920 41.060 ;
        RECT 168.165 40.340 168.915 40.510 ;
        RECT 162.870 39.600 163.390 40.140 ;
        RECT 163.560 39.770 165.210 40.290 ;
        RECT 165.380 39.600 167.070 40.120 ;
        RECT 162.180 38.510 163.390 39.600 ;
        RECT 163.560 38.510 167.070 39.600 ;
        RECT 168.165 39.520 168.515 40.170 ;
        RECT 168.685 39.350 168.915 40.340 ;
        RECT 168.165 39.180 168.915 39.350 ;
        RECT 168.165 38.680 168.420 39.180 ;
        RECT 168.590 38.510 168.920 39.010 ;
        RECT 169.090 38.680 169.260 40.800 ;
        RECT 169.620 40.700 169.950 41.060 ;
        RECT 170.120 40.670 170.615 40.840 ;
        RECT 170.820 40.670 171.675 40.840 ;
        RECT 169.490 39.480 169.950 40.530 ;
        RECT 169.430 38.695 169.755 39.480 ;
        RECT 170.120 39.310 170.290 40.670 ;
        RECT 170.460 39.760 170.810 40.380 ;
        RECT 170.980 40.160 171.335 40.380 ;
        RECT 170.980 39.570 171.150 40.160 ;
        RECT 171.505 39.960 171.675 40.670 ;
        RECT 172.550 40.600 172.880 41.060 ;
        RECT 173.090 40.700 173.440 40.870 ;
        RECT 171.880 40.130 172.670 40.380 ;
        RECT 173.090 40.310 173.350 40.700 ;
        RECT 173.660 40.610 174.610 40.890 ;
        RECT 174.780 40.620 174.970 41.060 ;
        RECT 175.140 40.680 176.210 40.850 ;
        RECT 172.840 39.960 173.010 40.140 ;
        RECT 170.120 39.140 170.515 39.310 ;
        RECT 170.685 39.180 171.150 39.570 ;
        RECT 171.320 39.790 173.010 39.960 ;
        RECT 170.345 39.010 170.515 39.140 ;
        RECT 171.320 39.010 171.490 39.790 ;
        RECT 173.180 39.620 173.350 40.310 ;
        RECT 171.850 39.450 173.350 39.620 ;
        RECT 173.540 39.650 173.750 40.440 ;
        RECT 173.920 39.820 174.270 40.440 ;
        RECT 174.440 39.830 174.610 40.610 ;
        RECT 175.140 40.450 175.310 40.680 ;
        RECT 174.780 40.280 175.310 40.450 ;
        RECT 174.780 40.000 175.000 40.280 ;
        RECT 175.480 40.110 175.720 40.510 ;
        RECT 174.440 39.660 174.845 39.830 ;
        RECT 175.180 39.740 175.720 40.110 ;
        RECT 175.890 40.325 176.210 40.680 ;
        RECT 176.455 40.600 176.760 41.060 ;
        RECT 176.930 40.350 177.185 40.880 ;
        RECT 175.890 40.150 176.215 40.325 ;
        RECT 175.890 39.850 176.805 40.150 ;
        RECT 176.065 39.820 176.805 39.850 ;
        RECT 173.540 39.490 174.215 39.650 ;
        RECT 174.675 39.570 174.845 39.660 ;
        RECT 173.540 39.480 174.505 39.490 ;
        RECT 173.180 39.310 173.350 39.450 ;
        RECT 169.925 38.510 170.175 38.970 ;
        RECT 170.345 38.680 170.595 39.010 ;
        RECT 170.810 38.680 171.490 39.010 ;
        RECT 171.660 39.110 172.735 39.280 ;
        RECT 173.180 39.140 173.740 39.310 ;
        RECT 174.045 39.190 174.505 39.480 ;
        RECT 174.675 39.400 175.895 39.570 ;
        RECT 171.660 38.770 171.830 39.110 ;
        RECT 172.065 38.510 172.395 38.940 ;
        RECT 172.565 38.770 172.735 39.110 ;
        RECT 173.030 38.510 173.400 38.970 ;
        RECT 173.570 38.680 173.740 39.140 ;
        RECT 174.675 39.020 174.845 39.400 ;
        RECT 176.065 39.230 176.235 39.820 ;
        RECT 176.975 39.700 177.185 40.350 ;
        RECT 173.975 38.680 174.845 39.020 ;
        RECT 175.435 39.060 176.235 39.230 ;
        RECT 175.015 38.510 175.265 38.970 ;
        RECT 175.435 38.770 175.605 39.060 ;
        RECT 175.785 38.510 176.115 38.890 ;
        RECT 176.455 38.510 176.760 39.650 ;
        RECT 176.930 38.820 177.185 39.700 ;
        RECT 177.365 40.320 177.620 40.890 ;
        RECT 177.790 40.660 178.120 41.060 ;
        RECT 178.545 40.525 179.075 40.890 ;
        RECT 179.265 40.720 179.540 40.890 ;
        RECT 179.260 40.550 179.540 40.720 ;
        RECT 178.545 40.490 178.720 40.525 ;
        RECT 177.790 40.320 178.720 40.490 ;
        RECT 177.365 39.650 177.535 40.320 ;
        RECT 177.790 40.150 177.960 40.320 ;
        RECT 177.705 39.820 177.960 40.150 ;
        RECT 178.185 39.820 178.380 40.150 ;
        RECT 177.365 38.680 177.700 39.650 ;
        RECT 177.870 38.510 178.040 39.650 ;
        RECT 178.210 38.850 178.380 39.820 ;
        RECT 178.550 39.190 178.720 40.320 ;
        RECT 178.890 39.530 179.060 40.330 ;
        RECT 179.265 39.730 179.540 40.550 ;
        RECT 179.710 39.530 179.900 40.890 ;
        RECT 180.080 40.525 180.590 41.060 ;
        RECT 180.810 40.250 181.055 40.855 ;
        RECT 181.500 40.290 183.170 41.060 ;
        RECT 183.805 40.320 184.060 40.890 ;
        RECT 184.230 40.660 184.560 41.060 ;
        RECT 184.985 40.525 185.515 40.890 ;
        RECT 185.705 40.720 185.980 40.890 ;
        RECT 185.700 40.550 185.980 40.720 ;
        RECT 184.985 40.490 185.160 40.525 ;
        RECT 184.230 40.320 185.160 40.490 ;
        RECT 180.100 40.080 181.330 40.250 ;
        RECT 178.890 39.360 179.900 39.530 ;
        RECT 180.070 39.515 180.820 39.705 ;
        RECT 178.550 39.020 179.675 39.190 ;
        RECT 180.070 38.850 180.240 39.515 ;
        RECT 180.990 39.270 181.330 40.080 ;
        RECT 181.500 39.770 182.250 40.290 ;
        RECT 182.420 39.600 183.170 40.120 ;
        RECT 178.210 38.680 180.240 38.850 ;
        RECT 180.410 38.510 180.580 39.270 ;
        RECT 180.815 38.860 181.330 39.270 ;
        RECT 181.500 38.510 183.170 39.600 ;
        RECT 183.805 39.650 183.975 40.320 ;
        RECT 184.230 40.150 184.400 40.320 ;
        RECT 184.145 39.820 184.400 40.150 ;
        RECT 184.625 39.820 184.820 40.150 ;
        RECT 183.805 38.680 184.140 39.650 ;
        RECT 184.310 38.510 184.480 39.650 ;
        RECT 184.650 38.850 184.820 39.820 ;
        RECT 184.990 39.190 185.160 40.320 ;
        RECT 185.330 39.530 185.500 40.330 ;
        RECT 185.705 39.730 185.980 40.550 ;
        RECT 186.150 39.530 186.340 40.890 ;
        RECT 186.520 40.525 187.030 41.060 ;
        RECT 187.250 40.250 187.495 40.855 ;
        RECT 187.940 40.335 188.230 41.060 ;
        RECT 188.400 40.310 189.610 41.060 ;
        RECT 189.785 40.320 190.040 40.890 ;
        RECT 190.210 40.660 190.540 41.060 ;
        RECT 190.965 40.525 191.495 40.890 ;
        RECT 190.965 40.490 191.140 40.525 ;
        RECT 190.210 40.320 191.140 40.490 ;
        RECT 191.685 40.380 191.960 40.890 ;
        RECT 186.540 40.080 187.770 40.250 ;
        RECT 185.330 39.360 186.340 39.530 ;
        RECT 186.510 39.515 187.260 39.705 ;
        RECT 184.990 39.020 186.115 39.190 ;
        RECT 186.510 38.850 186.680 39.515 ;
        RECT 187.430 39.270 187.770 40.080 ;
        RECT 188.400 39.770 188.920 40.310 ;
        RECT 184.650 38.680 186.680 38.850 ;
        RECT 186.850 38.510 187.020 39.270 ;
        RECT 187.255 38.860 187.770 39.270 ;
        RECT 187.940 38.510 188.230 39.675 ;
        RECT 189.090 39.600 189.610 40.140 ;
        RECT 188.400 38.510 189.610 39.600 ;
        RECT 189.785 39.650 189.955 40.320 ;
        RECT 190.210 40.150 190.380 40.320 ;
        RECT 190.125 39.820 190.380 40.150 ;
        RECT 190.605 39.820 190.800 40.150 ;
        RECT 189.785 38.680 190.120 39.650 ;
        RECT 190.290 38.510 190.460 39.650 ;
        RECT 190.630 38.850 190.800 39.820 ;
        RECT 190.970 39.190 191.140 40.320 ;
        RECT 191.310 39.530 191.480 40.330 ;
        RECT 191.680 40.210 191.960 40.380 ;
        RECT 191.685 39.730 191.960 40.210 ;
        RECT 192.130 39.530 192.320 40.890 ;
        RECT 192.500 40.525 193.010 41.060 ;
        RECT 193.230 40.250 193.475 40.855 ;
        RECT 193.920 40.310 195.130 41.060 ;
        RECT 195.305 40.510 195.560 40.800 ;
        RECT 195.730 40.680 196.060 41.060 ;
        RECT 195.305 40.340 196.055 40.510 ;
        RECT 192.520 40.080 193.750 40.250 ;
        RECT 191.310 39.360 192.320 39.530 ;
        RECT 192.490 39.515 193.240 39.705 ;
        RECT 190.970 39.020 192.095 39.190 ;
        RECT 192.490 38.850 192.660 39.515 ;
        RECT 193.410 39.270 193.750 40.080 ;
        RECT 193.920 39.770 194.440 40.310 ;
        RECT 194.610 39.600 195.130 40.140 ;
        RECT 190.630 38.680 192.660 38.850 ;
        RECT 192.830 38.510 193.000 39.270 ;
        RECT 193.235 38.860 193.750 39.270 ;
        RECT 193.920 38.510 195.130 39.600 ;
        RECT 195.305 39.520 195.655 40.170 ;
        RECT 195.825 39.350 196.055 40.340 ;
        RECT 195.305 39.180 196.055 39.350 ;
        RECT 195.305 38.680 195.560 39.180 ;
        RECT 195.730 38.510 196.060 39.010 ;
        RECT 196.230 38.680 196.400 40.800 ;
        RECT 196.760 40.700 197.090 41.060 ;
        RECT 197.260 40.670 197.755 40.840 ;
        RECT 197.960 40.670 198.815 40.840 ;
        RECT 196.630 39.480 197.090 40.530 ;
        RECT 196.570 38.695 196.895 39.480 ;
        RECT 197.260 39.310 197.430 40.670 ;
        RECT 197.600 39.760 197.950 40.380 ;
        RECT 198.120 40.160 198.475 40.380 ;
        RECT 198.120 39.570 198.290 40.160 ;
        RECT 198.645 39.960 198.815 40.670 ;
        RECT 199.690 40.600 200.020 41.060 ;
        RECT 200.230 40.700 200.580 40.870 ;
        RECT 199.020 40.130 199.810 40.380 ;
        RECT 200.230 40.310 200.490 40.700 ;
        RECT 200.800 40.610 201.750 40.890 ;
        RECT 201.920 40.620 202.110 41.060 ;
        RECT 202.280 40.680 203.350 40.850 ;
        RECT 199.980 39.960 200.150 40.140 ;
        RECT 197.260 39.140 197.655 39.310 ;
        RECT 197.825 39.180 198.290 39.570 ;
        RECT 198.460 39.790 200.150 39.960 ;
        RECT 197.485 39.010 197.655 39.140 ;
        RECT 198.460 39.010 198.630 39.790 ;
        RECT 200.320 39.620 200.490 40.310 ;
        RECT 198.990 39.450 200.490 39.620 ;
        RECT 200.680 39.650 200.890 40.440 ;
        RECT 201.060 39.820 201.410 40.440 ;
        RECT 201.580 39.830 201.750 40.610 ;
        RECT 202.280 40.450 202.450 40.680 ;
        RECT 201.920 40.280 202.450 40.450 ;
        RECT 201.920 40.000 202.140 40.280 ;
        RECT 202.620 40.110 202.860 40.510 ;
        RECT 201.580 39.660 201.985 39.830 ;
        RECT 202.320 39.740 202.860 40.110 ;
        RECT 203.030 40.325 203.350 40.680 ;
        RECT 203.595 40.600 203.900 41.060 ;
        RECT 204.070 40.350 204.325 40.880 ;
        RECT 203.030 40.150 203.355 40.325 ;
        RECT 203.030 39.850 203.945 40.150 ;
        RECT 203.205 39.820 203.945 39.850 ;
        RECT 200.680 39.490 201.355 39.650 ;
        RECT 201.815 39.570 201.985 39.660 ;
        RECT 200.680 39.480 201.645 39.490 ;
        RECT 200.320 39.310 200.490 39.450 ;
        RECT 197.065 38.510 197.315 38.970 ;
        RECT 197.485 38.680 197.735 39.010 ;
        RECT 197.950 38.680 198.630 39.010 ;
        RECT 198.800 39.110 199.875 39.280 ;
        RECT 200.320 39.140 200.880 39.310 ;
        RECT 201.185 39.190 201.645 39.480 ;
        RECT 201.815 39.400 203.035 39.570 ;
        RECT 198.800 38.770 198.970 39.110 ;
        RECT 199.205 38.510 199.535 38.940 ;
        RECT 199.705 38.770 199.875 39.110 ;
        RECT 200.170 38.510 200.540 38.970 ;
        RECT 200.710 38.680 200.880 39.140 ;
        RECT 201.815 39.020 201.985 39.400 ;
        RECT 203.205 39.230 203.375 39.820 ;
        RECT 204.115 39.700 204.325 40.350 ;
        RECT 201.115 38.680 201.985 39.020 ;
        RECT 202.575 39.060 203.375 39.230 ;
        RECT 202.155 38.510 202.405 38.970 ;
        RECT 202.575 38.770 202.745 39.060 ;
        RECT 202.925 38.510 203.255 38.890 ;
        RECT 203.595 38.510 203.900 39.650 ;
        RECT 204.070 38.820 204.325 39.700 ;
        RECT 204.505 40.320 204.760 40.890 ;
        RECT 204.930 40.660 205.260 41.060 ;
        RECT 205.685 40.525 206.215 40.890 ;
        RECT 206.405 40.720 206.680 40.890 ;
        RECT 206.400 40.550 206.680 40.720 ;
        RECT 205.685 40.490 205.860 40.525 ;
        RECT 204.930 40.320 205.860 40.490 ;
        RECT 204.505 39.650 204.675 40.320 ;
        RECT 204.930 40.150 205.100 40.320 ;
        RECT 204.845 39.820 205.100 40.150 ;
        RECT 205.325 39.820 205.520 40.150 ;
        RECT 204.505 38.680 204.840 39.650 ;
        RECT 205.010 38.510 205.180 39.650 ;
        RECT 205.350 38.850 205.520 39.820 ;
        RECT 205.690 39.190 205.860 40.320 ;
        RECT 206.030 39.530 206.200 40.330 ;
        RECT 206.405 39.730 206.680 40.550 ;
        RECT 206.850 39.530 207.040 40.890 ;
        RECT 207.220 40.525 207.730 41.060 ;
        RECT 207.950 40.250 208.195 40.855 ;
        RECT 208.640 40.310 209.850 41.060 ;
        RECT 210.135 40.430 210.420 40.890 ;
        RECT 210.590 40.600 210.860 41.060 ;
        RECT 207.240 40.080 208.470 40.250 ;
        RECT 206.030 39.360 207.040 39.530 ;
        RECT 207.210 39.515 207.960 39.705 ;
        RECT 205.690 39.020 206.815 39.190 ;
        RECT 207.210 38.850 207.380 39.515 ;
        RECT 208.130 39.270 208.470 40.080 ;
        RECT 208.640 39.770 209.160 40.310 ;
        RECT 210.135 40.260 211.090 40.430 ;
        RECT 209.330 39.600 209.850 40.140 ;
        RECT 205.350 38.680 207.380 38.850 ;
        RECT 207.550 38.510 207.720 39.270 ;
        RECT 207.955 38.860 208.470 39.270 ;
        RECT 208.640 38.510 209.850 39.600 ;
        RECT 210.020 39.530 210.710 40.090 ;
        RECT 210.880 39.360 211.090 40.260 ;
        RECT 210.135 39.140 211.090 39.360 ;
        RECT 211.260 40.090 211.660 40.890 ;
        RECT 211.850 40.430 212.130 40.890 ;
        RECT 212.650 40.600 212.975 41.060 ;
        RECT 211.850 40.260 212.975 40.430 ;
        RECT 213.145 40.320 213.530 40.890 ;
        RECT 213.700 40.335 213.990 41.060 ;
        RECT 214.165 40.510 214.420 40.800 ;
        RECT 214.590 40.680 214.920 41.060 ;
        RECT 214.165 40.340 214.915 40.510 ;
        RECT 212.525 40.150 212.975 40.260 ;
        RECT 211.260 39.530 212.355 40.090 ;
        RECT 212.525 39.820 213.080 40.150 ;
        RECT 210.135 38.680 210.420 39.140 ;
        RECT 210.590 38.510 210.860 38.970 ;
        RECT 211.260 38.680 211.660 39.530 ;
        RECT 212.525 39.360 212.975 39.820 ;
        RECT 213.250 39.650 213.530 40.320 ;
        RECT 211.850 39.140 212.975 39.360 ;
        RECT 211.850 38.680 212.130 39.140 ;
        RECT 212.650 38.510 212.975 38.970 ;
        RECT 213.145 38.680 213.530 39.650 ;
        RECT 213.700 38.510 213.990 39.675 ;
        RECT 214.165 39.520 214.515 40.170 ;
        RECT 214.685 39.350 214.915 40.340 ;
        RECT 214.165 39.180 214.915 39.350 ;
        RECT 214.165 38.680 214.420 39.180 ;
        RECT 214.590 38.510 214.920 39.010 ;
        RECT 215.090 38.680 215.260 40.800 ;
        RECT 215.620 40.700 215.950 41.060 ;
        RECT 216.120 40.670 216.615 40.840 ;
        RECT 216.820 40.670 217.675 40.840 ;
        RECT 215.490 39.480 215.950 40.530 ;
        RECT 215.430 38.695 215.755 39.480 ;
        RECT 216.120 39.310 216.290 40.670 ;
        RECT 216.460 39.760 216.810 40.380 ;
        RECT 216.980 40.160 217.335 40.380 ;
        RECT 216.980 39.570 217.150 40.160 ;
        RECT 217.505 39.960 217.675 40.670 ;
        RECT 218.550 40.600 218.880 41.060 ;
        RECT 219.090 40.700 219.440 40.870 ;
        RECT 217.880 40.130 218.670 40.380 ;
        RECT 219.090 40.310 219.350 40.700 ;
        RECT 219.660 40.610 220.610 40.890 ;
        RECT 220.780 40.620 220.970 41.060 ;
        RECT 221.140 40.680 222.210 40.850 ;
        RECT 218.840 39.960 219.010 40.140 ;
        RECT 216.120 39.140 216.515 39.310 ;
        RECT 216.685 39.180 217.150 39.570 ;
        RECT 217.320 39.790 219.010 39.960 ;
        RECT 216.345 39.010 216.515 39.140 ;
        RECT 217.320 39.010 217.490 39.790 ;
        RECT 219.180 39.620 219.350 40.310 ;
        RECT 217.850 39.450 219.350 39.620 ;
        RECT 219.540 39.650 219.750 40.440 ;
        RECT 219.920 39.820 220.270 40.440 ;
        RECT 220.440 39.830 220.610 40.610 ;
        RECT 221.140 40.450 221.310 40.680 ;
        RECT 220.780 40.280 221.310 40.450 ;
        RECT 220.780 40.000 221.000 40.280 ;
        RECT 221.480 40.110 221.720 40.510 ;
        RECT 220.440 39.660 220.845 39.830 ;
        RECT 221.180 39.740 221.720 40.110 ;
        RECT 221.890 40.325 222.210 40.680 ;
        RECT 222.455 40.600 222.760 41.060 ;
        RECT 222.930 40.350 223.185 40.880 ;
        RECT 221.890 40.150 222.215 40.325 ;
        RECT 221.890 39.850 222.805 40.150 ;
        RECT 222.065 39.820 222.805 39.850 ;
        RECT 219.540 39.490 220.215 39.650 ;
        RECT 220.675 39.570 220.845 39.660 ;
        RECT 219.540 39.480 220.505 39.490 ;
        RECT 219.180 39.310 219.350 39.450 ;
        RECT 215.925 38.510 216.175 38.970 ;
        RECT 216.345 38.680 216.595 39.010 ;
        RECT 216.810 38.680 217.490 39.010 ;
        RECT 217.660 39.110 218.735 39.280 ;
        RECT 219.180 39.140 219.740 39.310 ;
        RECT 220.045 39.190 220.505 39.480 ;
        RECT 220.675 39.400 221.895 39.570 ;
        RECT 217.660 38.770 217.830 39.110 ;
        RECT 218.065 38.510 218.395 38.940 ;
        RECT 218.565 38.770 218.735 39.110 ;
        RECT 219.030 38.510 219.400 38.970 ;
        RECT 219.570 38.680 219.740 39.140 ;
        RECT 220.675 39.020 220.845 39.400 ;
        RECT 222.065 39.230 222.235 39.820 ;
        RECT 222.975 39.700 223.185 40.350 ;
        RECT 219.975 38.680 220.845 39.020 ;
        RECT 221.435 39.060 222.235 39.230 ;
        RECT 221.015 38.510 221.265 38.970 ;
        RECT 221.435 38.770 221.605 39.060 ;
        RECT 221.785 38.510 222.115 38.890 ;
        RECT 222.455 38.510 222.760 39.650 ;
        RECT 222.930 38.820 223.185 39.700 ;
        RECT 223.395 40.320 224.010 40.890 ;
        RECT 224.180 40.550 224.395 41.060 ;
        RECT 224.625 40.550 224.905 40.880 ;
        RECT 225.085 40.550 225.325 41.060 ;
        RECT 223.395 39.300 223.710 40.320 ;
        RECT 223.880 39.650 224.050 40.150 ;
        RECT 224.300 39.820 224.565 40.380 ;
        RECT 224.735 39.650 224.905 40.550 ;
        RECT 225.075 39.820 225.430 40.380 ;
        RECT 225.665 40.320 225.920 40.890 ;
        RECT 226.090 40.660 226.420 41.060 ;
        RECT 226.845 40.525 227.375 40.890 ;
        RECT 227.565 40.720 227.840 40.890 ;
        RECT 227.560 40.550 227.840 40.720 ;
        RECT 226.845 40.490 227.020 40.525 ;
        RECT 226.090 40.320 227.020 40.490 ;
        RECT 225.665 39.650 225.835 40.320 ;
        RECT 226.090 40.150 226.260 40.320 ;
        RECT 226.005 39.820 226.260 40.150 ;
        RECT 226.485 39.820 226.680 40.150 ;
        RECT 223.880 39.480 225.305 39.650 ;
        RECT 223.395 38.680 223.930 39.300 ;
        RECT 224.100 38.510 224.430 39.310 ;
        RECT 224.915 39.305 225.305 39.480 ;
        RECT 225.665 38.680 226.000 39.650 ;
        RECT 226.170 38.510 226.340 39.650 ;
        RECT 226.510 38.850 226.680 39.820 ;
        RECT 226.850 39.190 227.020 40.320 ;
        RECT 227.190 39.530 227.360 40.330 ;
        RECT 227.565 39.730 227.840 40.550 ;
        RECT 228.010 39.530 228.200 40.890 ;
        RECT 228.380 40.525 228.890 41.060 ;
        RECT 229.110 40.250 229.355 40.855 ;
        RECT 229.805 40.320 230.060 40.890 ;
        RECT 230.230 40.660 230.560 41.060 ;
        RECT 230.985 40.525 231.515 40.890 ;
        RECT 230.985 40.490 231.160 40.525 ;
        RECT 230.230 40.320 231.160 40.490 ;
        RECT 228.400 40.080 229.630 40.250 ;
        RECT 227.190 39.360 228.200 39.530 ;
        RECT 228.370 39.515 229.120 39.705 ;
        RECT 226.850 39.020 227.975 39.190 ;
        RECT 228.370 38.850 228.540 39.515 ;
        RECT 229.290 39.270 229.630 40.080 ;
        RECT 226.510 38.680 228.540 38.850 ;
        RECT 228.710 38.510 228.880 39.270 ;
        RECT 229.115 38.860 229.630 39.270 ;
        RECT 229.805 39.650 229.975 40.320 ;
        RECT 230.230 40.150 230.400 40.320 ;
        RECT 230.145 39.820 230.400 40.150 ;
        RECT 230.625 39.820 230.820 40.150 ;
        RECT 229.805 38.680 230.140 39.650 ;
        RECT 230.310 38.510 230.480 39.650 ;
        RECT 230.650 38.850 230.820 39.820 ;
        RECT 230.990 39.190 231.160 40.320 ;
        RECT 231.330 39.530 231.500 40.330 ;
        RECT 231.705 40.040 231.980 40.890 ;
        RECT 231.700 39.870 231.980 40.040 ;
        RECT 231.705 39.730 231.980 39.870 ;
        RECT 232.150 39.530 232.340 40.890 ;
        RECT 232.520 40.525 233.030 41.060 ;
        RECT 233.250 40.250 233.495 40.855 ;
        RECT 234.055 40.430 234.340 40.890 ;
        RECT 234.510 40.600 234.780 41.060 ;
        RECT 234.055 40.260 235.010 40.430 ;
        RECT 232.540 40.080 233.770 40.250 ;
        RECT 231.330 39.360 232.340 39.530 ;
        RECT 232.510 39.515 233.260 39.705 ;
        RECT 230.990 39.020 232.115 39.190 ;
        RECT 232.510 38.850 232.680 39.515 ;
        RECT 233.430 39.270 233.770 40.080 ;
        RECT 233.940 39.530 234.630 40.090 ;
        RECT 234.800 39.360 235.010 40.260 ;
        RECT 230.650 38.680 232.680 38.850 ;
        RECT 232.850 38.510 233.020 39.270 ;
        RECT 233.255 38.860 233.770 39.270 ;
        RECT 234.055 39.140 235.010 39.360 ;
        RECT 235.180 40.090 235.580 40.890 ;
        RECT 235.770 40.430 236.050 40.890 ;
        RECT 236.570 40.600 236.895 41.060 ;
        RECT 235.770 40.260 236.895 40.430 ;
        RECT 237.065 40.320 237.450 40.890 ;
        RECT 237.625 40.660 237.960 41.060 ;
        RECT 238.130 40.490 238.335 40.890 ;
        RECT 238.545 40.580 238.820 41.060 ;
        RECT 239.030 40.560 239.290 40.890 ;
        RECT 236.445 40.150 236.895 40.260 ;
        RECT 235.180 39.530 236.275 40.090 ;
        RECT 236.445 39.820 237.000 40.150 ;
        RECT 234.055 38.680 234.340 39.140 ;
        RECT 234.510 38.510 234.780 38.970 ;
        RECT 235.180 38.680 235.580 39.530 ;
        RECT 236.445 39.360 236.895 39.820 ;
        RECT 237.170 39.650 237.450 40.320 ;
        RECT 235.770 39.140 236.895 39.360 ;
        RECT 235.770 38.680 236.050 39.140 ;
        RECT 236.570 38.510 236.895 38.970 ;
        RECT 237.065 38.680 237.450 39.650 ;
        RECT 237.650 40.320 238.335 40.490 ;
        RECT 237.650 39.290 237.990 40.320 ;
        RECT 238.160 39.650 238.410 40.150 ;
        RECT 238.590 39.820 238.950 40.400 ;
        RECT 239.120 39.650 239.290 40.560 ;
        RECT 239.460 40.335 239.750 41.060 ;
        RECT 239.920 40.310 241.130 41.060 ;
        RECT 241.305 40.320 241.560 40.890 ;
        RECT 241.730 40.660 242.060 41.060 ;
        RECT 242.485 40.525 243.015 40.890 ;
        RECT 242.485 40.490 242.660 40.525 ;
        RECT 241.730 40.320 242.660 40.490 ;
        RECT 243.205 40.380 243.480 40.890 ;
        RECT 239.920 39.770 240.440 40.310 ;
        RECT 238.160 39.480 239.290 39.650 ;
        RECT 237.650 39.115 238.315 39.290 ;
        RECT 237.625 38.510 237.960 38.935 ;
        RECT 238.130 38.710 238.315 39.115 ;
        RECT 238.520 38.510 238.850 39.290 ;
        RECT 239.020 38.710 239.290 39.480 ;
        RECT 239.460 38.510 239.750 39.675 ;
        RECT 240.610 39.600 241.130 40.140 ;
        RECT 239.920 38.510 241.130 39.600 ;
        RECT 241.305 39.650 241.475 40.320 ;
        RECT 241.730 40.150 241.900 40.320 ;
        RECT 241.645 39.820 241.900 40.150 ;
        RECT 242.125 39.820 242.320 40.150 ;
        RECT 241.305 38.680 241.640 39.650 ;
        RECT 241.810 38.510 241.980 39.650 ;
        RECT 242.150 38.850 242.320 39.820 ;
        RECT 242.490 39.190 242.660 40.320 ;
        RECT 242.830 39.530 243.000 40.330 ;
        RECT 243.200 40.210 243.480 40.380 ;
        RECT 243.205 39.730 243.480 40.210 ;
        RECT 243.650 39.530 243.840 40.890 ;
        RECT 244.020 40.525 244.530 41.060 ;
        RECT 244.750 40.250 244.995 40.855 ;
        RECT 245.445 40.320 245.700 40.890 ;
        RECT 245.870 40.660 246.200 41.060 ;
        RECT 246.625 40.525 247.155 40.890 ;
        RECT 246.625 40.490 246.800 40.525 ;
        RECT 245.870 40.320 246.800 40.490 ;
        RECT 244.040 40.080 245.270 40.250 ;
        RECT 242.830 39.360 243.840 39.530 ;
        RECT 244.010 39.515 244.760 39.705 ;
        RECT 242.490 39.020 243.615 39.190 ;
        RECT 244.010 38.850 244.180 39.515 ;
        RECT 244.930 39.270 245.270 40.080 ;
        RECT 242.150 38.680 244.180 38.850 ;
        RECT 244.350 38.510 244.520 39.270 ;
        RECT 244.755 38.860 245.270 39.270 ;
        RECT 245.445 39.650 245.615 40.320 ;
        RECT 245.870 40.150 246.040 40.320 ;
        RECT 245.785 39.820 246.040 40.150 ;
        RECT 246.265 39.820 246.460 40.150 ;
        RECT 245.445 38.680 245.780 39.650 ;
        RECT 245.950 38.510 246.120 39.650 ;
        RECT 246.290 38.850 246.460 39.820 ;
        RECT 246.630 39.190 246.800 40.320 ;
        RECT 246.970 39.530 247.140 40.330 ;
        RECT 247.345 40.040 247.620 40.890 ;
        RECT 247.340 39.870 247.620 40.040 ;
        RECT 247.345 39.730 247.620 39.870 ;
        RECT 247.790 39.530 247.980 40.890 ;
        RECT 248.160 40.525 248.670 41.060 ;
        RECT 248.890 40.250 249.135 40.855 ;
        RECT 249.580 40.320 249.965 40.890 ;
        RECT 250.135 40.600 250.460 41.060 ;
        RECT 250.980 40.430 251.260 40.890 ;
        RECT 248.180 40.080 249.410 40.250 ;
        RECT 246.970 39.360 247.980 39.530 ;
        RECT 248.150 39.515 248.900 39.705 ;
        RECT 246.630 39.020 247.755 39.190 ;
        RECT 248.150 38.850 248.320 39.515 ;
        RECT 249.070 39.270 249.410 40.080 ;
        RECT 246.290 38.680 248.320 38.850 ;
        RECT 248.490 38.510 248.660 39.270 ;
        RECT 248.895 38.860 249.410 39.270 ;
        RECT 249.580 39.650 249.860 40.320 ;
        RECT 250.135 40.260 251.260 40.430 ;
        RECT 250.135 40.150 250.585 40.260 ;
        RECT 250.030 39.820 250.585 40.150 ;
        RECT 251.450 40.090 251.850 40.890 ;
        RECT 252.250 40.600 252.520 41.060 ;
        RECT 252.690 40.430 252.975 40.890 ;
        RECT 249.580 38.680 249.965 39.650 ;
        RECT 250.135 39.360 250.585 39.820 ;
        RECT 250.755 39.530 251.850 40.090 ;
        RECT 250.135 39.140 251.260 39.360 ;
        RECT 250.135 38.510 250.460 38.970 ;
        RECT 250.980 38.680 251.260 39.140 ;
        RECT 251.450 38.680 251.850 39.530 ;
        RECT 252.020 40.260 252.975 40.430 ;
        RECT 253.260 40.310 254.470 41.060 ;
        RECT 254.640 40.680 255.530 40.850 ;
        RECT 252.020 39.360 252.230 40.260 ;
        RECT 252.400 39.530 253.090 40.090 ;
        RECT 253.260 39.770 253.780 40.310 ;
        RECT 253.950 39.600 254.470 40.140 ;
        RECT 254.640 40.125 255.190 40.510 ;
        RECT 255.360 39.955 255.530 40.680 ;
        RECT 252.020 39.140 252.975 39.360 ;
        RECT 252.250 38.510 252.520 38.970 ;
        RECT 252.690 38.680 252.975 39.140 ;
        RECT 253.260 38.510 254.470 39.600 ;
        RECT 254.640 39.885 255.530 39.955 ;
        RECT 255.700 40.380 255.920 40.840 ;
        RECT 256.090 40.520 256.340 41.060 ;
        RECT 256.510 40.410 256.770 40.890 ;
        RECT 257.155 40.590 257.440 41.060 ;
        RECT 257.610 40.420 257.940 40.890 ;
        RECT 258.110 40.590 258.280 41.060 ;
        RECT 258.450 40.420 258.780 40.890 ;
        RECT 258.950 40.590 259.120 41.060 ;
        RECT 259.290 40.420 259.620 40.890 ;
        RECT 259.790 40.590 259.960 41.060 ;
        RECT 260.130 40.420 260.460 40.890 ;
        RECT 255.700 40.355 255.950 40.380 ;
        RECT 255.700 39.930 256.030 40.355 ;
        RECT 254.640 39.860 255.535 39.885 ;
        RECT 254.640 39.845 255.545 39.860 ;
        RECT 254.640 39.830 255.550 39.845 ;
        RECT 254.640 39.825 255.560 39.830 ;
        RECT 254.640 39.815 255.565 39.825 ;
        RECT 254.640 39.805 255.570 39.815 ;
        RECT 254.640 39.800 255.580 39.805 ;
        RECT 254.640 39.790 255.590 39.800 ;
        RECT 254.640 39.785 255.600 39.790 ;
        RECT 254.640 39.335 254.900 39.785 ;
        RECT 255.265 39.780 255.600 39.785 ;
        RECT 255.265 39.775 255.615 39.780 ;
        RECT 255.265 39.765 255.630 39.775 ;
        RECT 255.265 39.760 255.655 39.765 ;
        RECT 256.200 39.760 256.430 40.155 ;
        RECT 255.265 39.755 256.430 39.760 ;
        RECT 255.295 39.720 256.430 39.755 ;
        RECT 255.330 39.695 256.430 39.720 ;
        RECT 255.360 39.665 256.430 39.695 ;
        RECT 255.380 39.635 256.430 39.665 ;
        RECT 255.400 39.605 256.430 39.635 ;
        RECT 255.470 39.595 256.430 39.605 ;
        RECT 255.495 39.585 256.430 39.595 ;
        RECT 255.515 39.570 256.430 39.585 ;
        RECT 255.535 39.555 256.430 39.570 ;
        RECT 255.540 39.545 256.325 39.555 ;
        RECT 255.555 39.510 256.325 39.545 ;
        RECT 255.070 39.190 255.400 39.435 ;
        RECT 255.570 39.260 256.325 39.510 ;
        RECT 256.600 39.380 256.770 40.410 ;
        RECT 256.940 40.240 260.460 40.420 ;
        RECT 260.630 40.240 260.905 41.060 ;
        RECT 256.940 39.700 257.340 40.240 ;
        RECT 261.080 40.115 261.420 40.890 ;
        RECT 261.590 40.600 261.760 41.060 ;
        RECT 262.000 40.625 262.360 40.890 ;
        RECT 262.000 40.620 262.355 40.625 ;
        RECT 262.000 40.610 262.350 40.620 ;
        RECT 262.000 40.605 262.345 40.610 ;
        RECT 262.000 40.595 262.340 40.605 ;
        RECT 262.990 40.600 263.160 41.060 ;
        RECT 262.000 40.590 262.335 40.595 ;
        RECT 262.000 40.580 262.325 40.590 ;
        RECT 262.000 40.570 262.315 40.580 ;
        RECT 262.000 40.430 262.300 40.570 ;
        RECT 261.590 40.240 262.300 40.430 ;
        RECT 262.490 40.430 262.820 40.510 ;
        RECT 263.330 40.430 263.670 40.890 ;
        RECT 262.490 40.240 263.670 40.430 ;
        RECT 263.840 40.310 265.050 41.060 ;
        RECT 265.220 40.335 265.510 41.060 ;
        RECT 265.680 40.320 266.065 40.890 ;
        RECT 266.235 40.600 266.560 41.060 ;
        RECT 267.080 40.430 267.360 40.890 ;
        RECT 257.510 39.870 258.875 40.070 ;
        RECT 259.195 39.870 260.855 40.070 ;
        RECT 256.940 39.400 258.700 39.700 ;
        RECT 255.070 39.165 255.255 39.190 ;
        RECT 254.640 39.065 255.255 39.165 ;
        RECT 254.640 38.510 255.245 39.065 ;
        RECT 255.420 38.680 255.900 39.020 ;
        RECT 256.070 38.510 256.325 39.055 ;
        RECT 256.495 38.680 256.770 39.380 ;
        RECT 257.105 38.850 257.520 39.230 ;
        RECT 257.690 39.020 257.860 39.400 ;
        RECT 258.030 38.850 258.360 39.210 ;
        RECT 258.530 39.020 258.700 39.400 ;
        RECT 258.870 39.480 260.905 39.690 ;
        RECT 258.870 38.850 259.200 39.480 ;
        RECT 257.105 38.680 259.200 38.850 ;
        RECT 259.370 38.510 259.620 39.310 ;
        RECT 259.790 38.680 259.960 39.480 ;
        RECT 260.130 38.510 260.460 39.310 ;
        RECT 260.630 38.680 260.905 39.480 ;
        RECT 261.080 38.680 261.360 40.115 ;
        RECT 261.590 39.670 261.875 40.240 ;
        RECT 262.060 39.840 262.530 40.070 ;
        RECT 262.700 40.050 263.030 40.070 ;
        RECT 262.700 39.870 263.150 40.050 ;
        RECT 263.340 39.870 263.670 40.070 ;
        RECT 261.590 39.455 262.740 39.670 ;
        RECT 261.530 38.510 262.240 39.285 ;
        RECT 262.410 38.680 262.740 39.455 ;
        RECT 262.935 38.755 263.150 39.870 ;
        RECT 263.440 39.530 263.670 39.870 ;
        RECT 263.840 39.770 264.360 40.310 ;
        RECT 264.530 39.600 265.050 40.140 ;
        RECT 263.330 38.510 263.660 39.230 ;
        RECT 263.840 38.510 265.050 39.600 ;
        RECT 265.220 38.510 265.510 39.675 ;
        RECT 265.680 39.650 265.960 40.320 ;
        RECT 266.235 40.260 267.360 40.430 ;
        RECT 266.235 40.150 266.685 40.260 ;
        RECT 266.130 39.820 266.685 40.150 ;
        RECT 267.550 40.090 267.950 40.890 ;
        RECT 268.350 40.600 268.620 41.060 ;
        RECT 268.790 40.430 269.075 40.890 ;
        RECT 265.680 38.680 266.065 39.650 ;
        RECT 266.235 39.360 266.685 39.820 ;
        RECT 266.855 39.530 267.950 40.090 ;
        RECT 266.235 39.140 267.360 39.360 ;
        RECT 266.235 38.510 266.560 38.970 ;
        RECT 267.080 38.680 267.360 39.140 ;
        RECT 267.550 38.680 267.950 39.530 ;
        RECT 268.120 40.260 269.075 40.430 ;
        RECT 268.120 39.360 268.330 40.260 ;
        RECT 270.340 40.240 270.550 41.060 ;
        RECT 270.720 40.260 271.050 40.890 ;
        RECT 268.500 39.530 269.190 40.090 ;
        RECT 270.720 39.660 270.970 40.260 ;
        RECT 271.220 40.240 271.450 41.060 ;
        RECT 271.660 40.410 271.920 40.855 ;
        RECT 272.195 40.580 272.365 41.060 ;
        RECT 272.575 40.410 272.905 40.860 ;
        RECT 273.075 40.580 273.245 41.060 ;
        RECT 273.430 40.560 273.665 40.890 ;
        RECT 273.835 40.660 274.165 41.060 ;
        RECT 273.430 40.410 273.600 40.560 ;
        RECT 274.335 40.490 274.505 40.840 ;
        RECT 274.675 40.660 275.065 41.060 ;
        RECT 275.235 40.540 275.490 40.840 ;
        RECT 275.870 40.660 276.200 41.060 ;
        RECT 275.235 40.490 275.630 40.540 ;
        RECT 276.370 40.490 276.540 40.760 ;
        RECT 276.710 40.660 277.040 41.060 ;
        RECT 277.210 40.490 277.465 40.760 ;
        RECT 273.825 40.425 275.630 40.490 ;
        RECT 271.660 40.240 272.340 40.410 ;
        RECT 271.140 39.820 271.470 40.070 ;
        RECT 268.120 39.140 269.075 39.360 ;
        RECT 268.350 38.510 268.620 38.970 ;
        RECT 268.790 38.680 269.075 39.140 ;
        RECT 270.340 38.510 270.550 39.650 ;
        RECT 270.720 38.680 271.050 39.660 ;
        RECT 271.220 38.510 271.450 39.650 ;
        RECT 271.660 39.505 272.000 40.070 ;
        RECT 272.170 39.335 272.340 40.240 ;
        RECT 272.510 40.240 273.600 40.410 ;
        RECT 273.770 40.320 275.630 40.425 ;
        RECT 273.770 40.255 273.975 40.320 ;
        RECT 272.510 39.730 272.680 40.240 ;
        RECT 273.770 40.070 273.940 40.255 ;
        RECT 272.850 39.900 273.940 40.070 ;
        RECT 274.110 39.730 274.295 40.150 ;
        RECT 272.510 39.445 273.795 39.730 ;
        RECT 273.975 39.445 274.295 39.730 ;
        RECT 274.465 39.445 274.775 40.150 ;
        RECT 274.965 39.820 275.255 40.150 ;
        RECT 271.660 39.275 272.340 39.335 ;
        RECT 274.965 39.275 275.195 39.820 ;
        RECT 271.660 39.105 275.195 39.275 ;
        RECT 271.660 38.925 271.920 39.105 ;
        RECT 275.425 38.935 275.630 40.320 ;
        RECT 275.800 39.480 276.070 40.490 ;
        RECT 276.240 40.320 277.465 40.490 ;
        RECT 277.650 40.330 277.950 41.060 ;
        RECT 276.240 39.650 276.410 40.320 ;
        RECT 278.130 40.150 278.360 40.770 ;
        RECT 278.560 40.500 278.785 40.880 ;
        RECT 278.955 40.670 279.285 41.060 ;
        RECT 278.560 40.320 278.890 40.500 ;
        RECT 276.580 39.820 276.960 40.150 ;
        RECT 277.130 39.820 277.465 40.150 ;
        RECT 277.655 39.820 277.950 40.150 ;
        RECT 278.130 39.820 278.545 40.150 ;
        RECT 276.240 39.480 276.555 39.650 ;
        RECT 272.125 38.510 272.485 38.935 ;
        RECT 272.995 38.510 273.325 38.935 ;
        RECT 273.830 38.510 274.170 38.935 ;
        RECT 275.095 38.720 275.630 38.935 ;
        RECT 275.805 38.510 276.120 39.310 ;
        RECT 276.385 39.020 276.555 39.480 ;
        RECT 276.725 39.140 276.960 39.820 ;
        RECT 278.715 39.650 278.890 40.320 ;
        RECT 279.060 39.820 279.300 40.470 ;
        RECT 279.940 40.320 280.325 40.890 ;
        RECT 280.495 40.600 280.820 41.060 ;
        RECT 281.340 40.430 281.620 40.890 ;
        RECT 279.940 39.650 280.220 40.320 ;
        RECT 280.495 40.260 281.620 40.430 ;
        RECT 280.495 40.150 280.945 40.260 ;
        RECT 280.390 39.820 280.945 40.150 ;
        RECT 281.810 40.090 282.210 40.890 ;
        RECT 282.610 40.600 282.880 41.060 ;
        RECT 283.050 40.430 283.335 40.890 ;
        RECT 283.620 40.515 288.965 41.060 ;
        RECT 276.320 38.865 276.555 39.020 ;
        RECT 277.130 38.865 277.465 39.650 ;
        RECT 276.320 38.850 277.465 38.865 ;
        RECT 276.385 38.695 277.465 38.850 ;
        RECT 277.650 39.290 278.545 39.620 ;
        RECT 278.715 39.460 279.300 39.650 ;
        RECT 277.650 39.120 278.855 39.290 ;
        RECT 277.650 38.690 277.980 39.120 ;
        RECT 278.160 38.510 278.355 38.950 ;
        RECT 278.525 38.690 278.855 39.120 ;
        RECT 279.025 38.690 279.300 39.460 ;
        RECT 279.940 38.680 280.325 39.650 ;
        RECT 280.495 39.360 280.945 39.820 ;
        RECT 281.115 39.530 282.210 40.090 ;
        RECT 280.495 39.140 281.620 39.360 ;
        RECT 280.495 38.510 280.820 38.970 ;
        RECT 281.340 38.680 281.620 39.140 ;
        RECT 281.810 38.680 282.210 39.530 ;
        RECT 282.380 40.260 283.335 40.430 ;
        RECT 282.380 39.360 282.590 40.260 ;
        RECT 282.760 39.530 283.450 40.090 ;
        RECT 285.205 39.685 285.545 40.515 ;
        RECT 289.140 40.290 290.810 41.060 ;
        RECT 290.980 40.335 291.270 41.060 ;
        RECT 291.440 40.515 296.785 41.060 ;
        RECT 282.380 39.140 283.335 39.360 ;
        RECT 282.610 38.510 282.880 38.970 ;
        RECT 283.050 38.680 283.335 39.140 ;
        RECT 287.025 38.945 287.375 40.195 ;
        RECT 289.140 39.770 289.890 40.290 ;
        RECT 290.060 39.600 290.810 40.120 ;
        RECT 293.025 39.685 293.365 40.515 ;
        RECT 296.960 40.290 299.550 41.060 ;
        RECT 299.725 40.350 299.980 40.880 ;
        RECT 300.150 40.600 300.455 41.060 ;
        RECT 300.700 40.680 301.770 40.850 ;
        RECT 283.620 38.510 288.965 38.945 ;
        RECT 289.140 38.510 290.810 39.600 ;
        RECT 290.980 38.510 291.270 39.675 ;
        RECT 294.845 38.945 295.195 40.195 ;
        RECT 296.960 39.770 298.170 40.290 ;
        RECT 298.340 39.600 299.550 40.120 ;
        RECT 291.440 38.510 296.785 38.945 ;
        RECT 296.960 38.510 299.550 39.600 ;
        RECT 299.725 39.700 299.935 40.350 ;
        RECT 300.700 40.325 301.020 40.680 ;
        RECT 300.695 40.150 301.020 40.325 ;
        RECT 300.105 39.850 301.020 40.150 ;
        RECT 301.190 40.110 301.430 40.510 ;
        RECT 301.600 40.450 301.770 40.680 ;
        RECT 301.940 40.620 302.130 41.060 ;
        RECT 302.300 40.610 303.250 40.890 ;
        RECT 303.470 40.700 303.820 40.870 ;
        RECT 301.600 40.280 302.130 40.450 ;
        RECT 300.105 39.820 300.845 39.850 ;
        RECT 299.725 38.820 299.980 39.700 ;
        RECT 300.150 38.510 300.455 39.650 ;
        RECT 300.675 39.230 300.845 39.820 ;
        RECT 301.190 39.740 301.730 40.110 ;
        RECT 301.910 40.000 302.130 40.280 ;
        RECT 302.300 39.830 302.470 40.610 ;
        RECT 302.065 39.660 302.470 39.830 ;
        RECT 302.640 39.820 302.990 40.440 ;
        RECT 302.065 39.570 302.235 39.660 ;
        RECT 303.160 39.650 303.370 40.440 ;
        RECT 301.015 39.400 302.235 39.570 ;
        RECT 302.695 39.490 303.370 39.650 ;
        RECT 300.675 39.060 301.475 39.230 ;
        RECT 300.795 38.510 301.125 38.890 ;
        RECT 301.305 38.770 301.475 39.060 ;
        RECT 302.065 39.020 302.235 39.400 ;
        RECT 302.405 39.480 303.370 39.490 ;
        RECT 303.560 40.310 303.820 40.700 ;
        RECT 304.030 40.600 304.360 41.060 ;
        RECT 305.235 40.670 306.090 40.840 ;
        RECT 306.295 40.670 306.790 40.840 ;
        RECT 306.960 40.700 307.290 41.060 ;
        RECT 303.560 39.620 303.730 40.310 ;
        RECT 303.900 39.960 304.070 40.140 ;
        RECT 304.240 40.130 305.030 40.380 ;
        RECT 305.235 39.960 305.405 40.670 ;
        RECT 305.575 40.160 305.930 40.380 ;
        RECT 303.900 39.790 305.590 39.960 ;
        RECT 302.405 39.190 302.865 39.480 ;
        RECT 303.560 39.450 305.060 39.620 ;
        RECT 303.560 39.310 303.730 39.450 ;
        RECT 303.170 39.140 303.730 39.310 ;
        RECT 301.645 38.510 301.895 38.970 ;
        RECT 302.065 38.680 302.935 39.020 ;
        RECT 303.170 38.680 303.340 39.140 ;
        RECT 304.175 39.110 305.250 39.280 ;
        RECT 303.510 38.510 303.880 38.970 ;
        RECT 304.175 38.770 304.345 39.110 ;
        RECT 304.515 38.510 304.845 38.940 ;
        RECT 305.080 38.770 305.250 39.110 ;
        RECT 305.420 39.010 305.590 39.790 ;
        RECT 305.760 39.570 305.930 40.160 ;
        RECT 306.100 39.760 306.450 40.380 ;
        RECT 305.760 39.180 306.225 39.570 ;
        RECT 306.620 39.310 306.790 40.670 ;
        RECT 306.960 39.480 307.420 40.530 ;
        RECT 306.395 39.140 306.790 39.310 ;
        RECT 306.395 39.010 306.565 39.140 ;
        RECT 305.420 38.680 306.100 39.010 ;
        RECT 306.315 38.680 306.565 39.010 ;
        RECT 306.735 38.510 306.985 38.970 ;
        RECT 307.155 38.695 307.480 39.480 ;
        RECT 307.650 38.680 307.820 40.800 ;
        RECT 307.990 40.680 308.320 41.060 ;
        RECT 308.490 40.510 308.745 40.800 ;
        RECT 307.995 40.340 308.745 40.510 ;
        RECT 307.995 39.350 308.225 40.340 ;
        RECT 309.840 40.310 311.050 41.060 ;
        RECT 308.395 39.520 308.745 40.170 ;
        RECT 309.840 39.600 310.360 40.140 ;
        RECT 310.530 39.770 311.050 40.310 ;
        RECT 307.995 39.180 308.745 39.350 ;
        RECT 307.990 38.510 308.320 39.010 ;
        RECT 308.490 38.680 308.745 39.180 ;
        RECT 309.840 38.510 311.050 39.600 ;
        RECT 162.095 38.340 311.135 38.510 ;
        RECT 162.180 37.250 163.390 38.340 ;
        RECT 163.560 37.250 167.070 38.340 ;
        RECT 162.180 36.540 162.700 37.080 ;
        RECT 162.870 36.710 163.390 37.250 ;
        RECT 163.560 36.560 165.210 37.080 ;
        RECT 165.380 36.730 167.070 37.250 ;
        RECT 167.240 37.200 167.625 38.170 ;
        RECT 167.795 37.880 168.120 38.340 ;
        RECT 168.640 37.710 168.920 38.170 ;
        RECT 167.795 37.490 168.920 37.710 ;
        RECT 162.180 35.790 163.390 36.540 ;
        RECT 163.560 35.790 167.070 36.560 ;
        RECT 167.240 36.530 167.520 37.200 ;
        RECT 167.795 37.030 168.245 37.490 ;
        RECT 169.110 37.320 169.510 38.170 ;
        RECT 169.910 37.880 170.180 38.340 ;
        RECT 170.350 37.710 170.635 38.170 ;
        RECT 167.690 36.700 168.245 37.030 ;
        RECT 168.415 36.760 169.510 37.320 ;
        RECT 167.795 36.590 168.245 36.700 ;
        RECT 167.240 35.960 167.625 36.530 ;
        RECT 167.795 36.420 168.920 36.590 ;
        RECT 167.795 35.790 168.120 36.250 ;
        RECT 168.640 35.960 168.920 36.420 ;
        RECT 169.110 35.960 169.510 36.760 ;
        RECT 169.680 37.490 170.635 37.710 ;
        RECT 169.680 36.590 169.890 37.490 ;
        RECT 170.060 36.760 170.750 37.320 ;
        RECT 170.925 37.200 171.260 38.170 ;
        RECT 171.430 37.200 171.600 38.340 ;
        RECT 171.770 38.000 173.800 38.170 ;
        RECT 169.680 36.420 170.635 36.590 ;
        RECT 169.910 35.790 170.180 36.250 ;
        RECT 170.350 35.960 170.635 36.420 ;
        RECT 170.925 36.530 171.095 37.200 ;
        RECT 171.770 37.030 171.940 38.000 ;
        RECT 171.265 36.700 171.520 37.030 ;
        RECT 171.745 36.700 171.940 37.030 ;
        RECT 172.110 37.660 173.235 37.830 ;
        RECT 171.350 36.530 171.520 36.700 ;
        RECT 172.110 36.530 172.280 37.660 ;
        RECT 170.925 35.960 171.180 36.530 ;
        RECT 171.350 36.360 172.280 36.530 ;
        RECT 172.450 37.320 173.460 37.490 ;
        RECT 172.450 36.520 172.620 37.320 ;
        RECT 172.825 36.640 173.100 37.120 ;
        RECT 172.820 36.470 173.100 36.640 ;
        RECT 172.105 36.325 172.280 36.360 ;
        RECT 171.350 35.790 171.680 36.190 ;
        RECT 172.105 35.960 172.635 36.325 ;
        RECT 172.825 35.960 173.100 36.470 ;
        RECT 173.270 35.960 173.460 37.320 ;
        RECT 173.630 37.335 173.800 38.000 ;
        RECT 173.970 37.580 174.140 38.340 ;
        RECT 174.375 37.580 174.890 37.990 ;
        RECT 173.630 37.145 174.380 37.335 ;
        RECT 174.550 36.770 174.890 37.580 ;
        RECT 175.060 37.175 175.350 38.340 ;
        RECT 175.525 37.200 175.860 38.170 ;
        RECT 176.030 37.200 176.200 38.340 ;
        RECT 176.370 38.000 178.400 38.170 ;
        RECT 173.660 36.600 174.890 36.770 ;
        RECT 173.640 35.790 174.150 36.325 ;
        RECT 174.370 35.995 174.615 36.600 ;
        RECT 175.525 36.530 175.695 37.200 ;
        RECT 176.370 37.030 176.540 38.000 ;
        RECT 175.865 36.700 176.120 37.030 ;
        RECT 176.345 36.700 176.540 37.030 ;
        RECT 176.710 37.660 177.835 37.830 ;
        RECT 175.950 36.530 176.120 36.700 ;
        RECT 176.710 36.530 176.880 37.660 ;
        RECT 175.060 35.790 175.350 36.515 ;
        RECT 175.525 35.960 175.780 36.530 ;
        RECT 175.950 36.360 176.880 36.530 ;
        RECT 177.050 37.320 178.060 37.490 ;
        RECT 177.050 36.520 177.220 37.320 ;
        RECT 176.705 36.325 176.880 36.360 ;
        RECT 175.950 35.790 176.280 36.190 ;
        RECT 176.705 35.960 177.235 36.325 ;
        RECT 177.425 36.300 177.700 37.120 ;
        RECT 177.420 36.130 177.700 36.300 ;
        RECT 177.425 35.960 177.700 36.130 ;
        RECT 177.870 35.960 178.060 37.320 ;
        RECT 178.230 37.335 178.400 38.000 ;
        RECT 178.570 37.580 178.740 38.340 ;
        RECT 178.975 37.580 179.490 37.990 ;
        RECT 178.230 37.145 178.980 37.335 ;
        RECT 179.150 36.770 179.490 37.580 ;
        RECT 180.695 37.710 180.980 38.170 ;
        RECT 181.150 37.880 181.420 38.340 ;
        RECT 180.695 37.490 181.650 37.710 ;
        RECT 178.260 36.600 179.490 36.770 ;
        RECT 180.580 36.760 181.270 37.320 ;
        RECT 178.240 35.790 178.750 36.325 ;
        RECT 178.970 35.995 179.215 36.600 ;
        RECT 181.440 36.590 181.650 37.490 ;
        RECT 180.695 36.420 181.650 36.590 ;
        RECT 181.820 37.320 182.220 38.170 ;
        RECT 182.410 37.710 182.690 38.170 ;
        RECT 183.210 37.880 183.535 38.340 ;
        RECT 182.410 37.490 183.535 37.710 ;
        RECT 181.820 36.760 182.915 37.320 ;
        RECT 183.085 37.030 183.535 37.490 ;
        RECT 183.705 37.200 184.090 38.170 ;
        RECT 184.265 37.670 184.520 38.170 ;
        RECT 184.690 37.840 185.020 38.340 ;
        RECT 184.265 37.500 185.015 37.670 ;
        RECT 180.695 35.960 180.980 36.420 ;
        RECT 181.150 35.790 181.420 36.250 ;
        RECT 181.820 35.960 182.220 36.760 ;
        RECT 183.085 36.700 183.640 37.030 ;
        RECT 183.085 36.590 183.535 36.700 ;
        RECT 182.410 36.420 183.535 36.590 ;
        RECT 183.810 36.530 184.090 37.200 ;
        RECT 184.265 36.680 184.615 37.330 ;
        RECT 182.410 35.960 182.690 36.420 ;
        RECT 183.210 35.790 183.535 36.250 ;
        RECT 183.705 35.960 184.090 36.530 ;
        RECT 184.785 36.510 185.015 37.500 ;
        RECT 184.265 36.340 185.015 36.510 ;
        RECT 184.265 36.050 184.520 36.340 ;
        RECT 184.690 35.790 185.020 36.170 ;
        RECT 185.190 36.050 185.360 38.170 ;
        RECT 185.530 37.370 185.855 38.155 ;
        RECT 186.025 37.880 186.275 38.340 ;
        RECT 186.445 37.840 186.695 38.170 ;
        RECT 186.910 37.840 187.590 38.170 ;
        RECT 186.445 37.710 186.615 37.840 ;
        RECT 186.220 37.540 186.615 37.710 ;
        RECT 185.590 36.320 186.050 37.370 ;
        RECT 186.220 36.180 186.390 37.540 ;
        RECT 186.785 37.280 187.250 37.670 ;
        RECT 186.560 36.470 186.910 37.090 ;
        RECT 187.080 36.690 187.250 37.280 ;
        RECT 187.420 37.060 187.590 37.840 ;
        RECT 187.760 37.740 187.930 38.080 ;
        RECT 188.165 37.910 188.495 38.340 ;
        RECT 188.665 37.740 188.835 38.080 ;
        RECT 189.130 37.880 189.500 38.340 ;
        RECT 187.760 37.570 188.835 37.740 ;
        RECT 189.670 37.710 189.840 38.170 ;
        RECT 190.075 37.830 190.945 38.170 ;
        RECT 191.115 37.880 191.365 38.340 ;
        RECT 189.280 37.540 189.840 37.710 ;
        RECT 189.280 37.400 189.450 37.540 ;
        RECT 187.950 37.230 189.450 37.400 ;
        RECT 190.145 37.370 190.605 37.660 ;
        RECT 187.420 36.890 189.110 37.060 ;
        RECT 187.080 36.470 187.435 36.690 ;
        RECT 187.605 36.180 187.775 36.890 ;
        RECT 187.980 36.470 188.770 36.720 ;
        RECT 188.940 36.710 189.110 36.890 ;
        RECT 189.280 36.540 189.450 37.230 ;
        RECT 185.720 35.790 186.050 36.150 ;
        RECT 186.220 36.010 186.715 36.180 ;
        RECT 186.920 36.010 187.775 36.180 ;
        RECT 188.650 35.790 188.980 36.250 ;
        RECT 189.190 36.150 189.450 36.540 ;
        RECT 189.640 37.360 190.605 37.370 ;
        RECT 190.775 37.450 190.945 37.830 ;
        RECT 191.535 37.790 191.705 38.080 ;
        RECT 191.885 37.960 192.215 38.340 ;
        RECT 191.535 37.620 192.335 37.790 ;
        RECT 189.640 37.200 190.315 37.360 ;
        RECT 190.775 37.280 191.995 37.450 ;
        RECT 189.640 36.410 189.850 37.200 ;
        RECT 190.775 37.190 190.945 37.280 ;
        RECT 190.020 36.410 190.370 37.030 ;
        RECT 190.540 37.020 190.945 37.190 ;
        RECT 190.540 36.240 190.710 37.020 ;
        RECT 190.880 36.570 191.100 36.850 ;
        RECT 191.280 36.740 191.820 37.110 ;
        RECT 192.165 37.030 192.335 37.620 ;
        RECT 192.555 37.200 192.860 38.340 ;
        RECT 193.030 37.150 193.285 38.030 ;
        RECT 192.165 37.000 192.905 37.030 ;
        RECT 190.880 36.400 191.410 36.570 ;
        RECT 189.190 35.980 189.540 36.150 ;
        RECT 189.760 35.960 190.710 36.240 ;
        RECT 190.880 35.790 191.070 36.230 ;
        RECT 191.240 36.170 191.410 36.400 ;
        RECT 191.580 36.340 191.820 36.740 ;
        RECT 191.990 36.700 192.905 37.000 ;
        RECT 191.990 36.525 192.315 36.700 ;
        RECT 191.990 36.170 192.310 36.525 ;
        RECT 193.075 36.500 193.285 37.150 ;
        RECT 191.240 36.000 192.310 36.170 ;
        RECT 192.555 35.790 192.860 36.250 ;
        RECT 193.030 35.970 193.285 36.500 ;
        RECT 193.460 37.200 193.845 38.170 ;
        RECT 194.015 37.880 194.340 38.340 ;
        RECT 194.860 37.710 195.140 38.170 ;
        RECT 194.015 37.490 195.140 37.710 ;
        RECT 193.460 36.530 193.740 37.200 ;
        RECT 194.015 37.030 194.465 37.490 ;
        RECT 195.330 37.320 195.730 38.170 ;
        RECT 196.130 37.880 196.400 38.340 ;
        RECT 196.570 37.710 196.855 38.170 ;
        RECT 193.910 36.700 194.465 37.030 ;
        RECT 194.635 36.760 195.730 37.320 ;
        RECT 194.015 36.590 194.465 36.700 ;
        RECT 193.460 35.960 193.845 36.530 ;
        RECT 194.015 36.420 195.140 36.590 ;
        RECT 194.015 35.790 194.340 36.250 ;
        RECT 194.860 35.960 195.140 36.420 ;
        RECT 195.330 35.960 195.730 36.760 ;
        RECT 195.900 37.490 196.855 37.710 ;
        RECT 197.255 37.710 197.540 38.170 ;
        RECT 197.710 37.880 197.980 38.340 ;
        RECT 197.255 37.490 198.210 37.710 ;
        RECT 195.900 36.590 196.110 37.490 ;
        RECT 196.280 36.760 196.970 37.320 ;
        RECT 197.140 36.760 197.830 37.320 ;
        RECT 198.000 36.590 198.210 37.490 ;
        RECT 195.900 36.420 196.855 36.590 ;
        RECT 196.130 35.790 196.400 36.250 ;
        RECT 196.570 35.960 196.855 36.420 ;
        RECT 197.255 36.420 198.210 36.590 ;
        RECT 198.380 37.320 198.780 38.170 ;
        RECT 198.970 37.710 199.250 38.170 ;
        RECT 199.770 37.880 200.095 38.340 ;
        RECT 198.970 37.490 200.095 37.710 ;
        RECT 198.380 36.760 199.475 37.320 ;
        RECT 199.645 37.030 200.095 37.490 ;
        RECT 200.265 37.200 200.650 38.170 ;
        RECT 197.255 35.960 197.540 36.420 ;
        RECT 197.710 35.790 197.980 36.250 ;
        RECT 198.380 35.960 198.780 36.760 ;
        RECT 199.645 36.700 200.200 37.030 ;
        RECT 199.645 36.590 200.095 36.700 ;
        RECT 198.970 36.420 200.095 36.590 ;
        RECT 200.370 36.530 200.650 37.200 ;
        RECT 200.820 37.175 201.110 38.340 ;
        RECT 201.280 37.250 203.870 38.340 ;
        RECT 198.970 35.960 199.250 36.420 ;
        RECT 199.770 35.790 200.095 36.250 ;
        RECT 200.265 35.960 200.650 36.530 ;
        RECT 201.280 36.560 202.490 37.080 ;
        RECT 202.660 36.730 203.870 37.250 ;
        RECT 204.505 37.200 204.840 38.170 ;
        RECT 205.010 37.200 205.180 38.340 ;
        RECT 205.350 38.000 207.380 38.170 ;
        RECT 200.820 35.790 201.110 36.515 ;
        RECT 201.280 35.790 203.870 36.560 ;
        RECT 204.505 36.530 204.675 37.200 ;
        RECT 205.350 37.030 205.520 38.000 ;
        RECT 204.845 36.700 205.100 37.030 ;
        RECT 205.325 36.700 205.520 37.030 ;
        RECT 205.690 37.660 206.815 37.830 ;
        RECT 204.930 36.530 205.100 36.700 ;
        RECT 205.690 36.530 205.860 37.660 ;
        RECT 204.505 35.960 204.760 36.530 ;
        RECT 204.930 36.360 205.860 36.530 ;
        RECT 206.030 37.320 207.040 37.490 ;
        RECT 206.030 36.520 206.200 37.320 ;
        RECT 206.405 36.640 206.680 37.120 ;
        RECT 206.400 36.470 206.680 36.640 ;
        RECT 205.685 36.325 205.860 36.360 ;
        RECT 204.930 35.790 205.260 36.190 ;
        RECT 205.685 35.960 206.215 36.325 ;
        RECT 206.405 35.960 206.680 36.470 ;
        RECT 206.850 35.960 207.040 37.320 ;
        RECT 207.210 37.335 207.380 38.000 ;
        RECT 207.550 37.580 207.720 38.340 ;
        RECT 207.955 37.580 208.470 37.990 ;
        RECT 207.210 37.145 207.960 37.335 ;
        RECT 208.130 36.770 208.470 37.580 ;
        RECT 208.640 37.250 210.310 38.340 ;
        RECT 207.240 36.600 208.470 36.770 ;
        RECT 207.220 35.790 207.730 36.325 ;
        RECT 207.950 35.995 208.195 36.600 ;
        RECT 208.640 36.560 209.390 37.080 ;
        RECT 209.560 36.730 210.310 37.250 ;
        RECT 210.940 37.580 211.455 37.990 ;
        RECT 211.690 37.580 211.860 38.340 ;
        RECT 212.030 38.000 214.060 38.170 ;
        RECT 210.940 36.770 211.280 37.580 ;
        RECT 212.030 37.335 212.200 38.000 ;
        RECT 212.595 37.660 213.720 37.830 ;
        RECT 211.450 37.145 212.200 37.335 ;
        RECT 212.370 37.320 213.380 37.490 ;
        RECT 210.940 36.600 212.170 36.770 ;
        RECT 208.640 35.790 210.310 36.560 ;
        RECT 211.215 35.995 211.460 36.600 ;
        RECT 211.680 35.790 212.190 36.325 ;
        RECT 212.370 35.960 212.560 37.320 ;
        RECT 212.730 36.640 213.005 37.120 ;
        RECT 212.730 36.470 213.010 36.640 ;
        RECT 213.210 36.520 213.380 37.320 ;
        RECT 213.550 36.530 213.720 37.660 ;
        RECT 213.890 37.030 214.060 38.000 ;
        RECT 214.230 37.200 214.400 38.340 ;
        RECT 214.570 37.200 214.905 38.170 ;
        RECT 213.890 36.700 214.085 37.030 ;
        RECT 214.310 36.700 214.565 37.030 ;
        RECT 214.310 36.530 214.480 36.700 ;
        RECT 214.735 36.530 214.905 37.200 ;
        RECT 212.730 35.960 213.005 36.470 ;
        RECT 213.550 36.360 214.480 36.530 ;
        RECT 213.550 36.325 213.725 36.360 ;
        RECT 213.195 35.960 213.725 36.325 ;
        RECT 214.150 35.790 214.480 36.190 ;
        RECT 214.650 35.960 214.905 36.530 ;
        RECT 215.085 37.200 215.420 38.170 ;
        RECT 215.590 37.200 215.760 38.340 ;
        RECT 215.930 38.000 217.960 38.170 ;
        RECT 215.085 36.530 215.255 37.200 ;
        RECT 215.930 37.030 216.100 38.000 ;
        RECT 215.425 36.700 215.680 37.030 ;
        RECT 215.905 36.700 216.100 37.030 ;
        RECT 216.270 37.660 217.395 37.830 ;
        RECT 215.510 36.530 215.680 36.700 ;
        RECT 216.270 36.530 216.440 37.660 ;
        RECT 215.085 35.960 215.340 36.530 ;
        RECT 215.510 36.360 216.440 36.530 ;
        RECT 216.610 37.320 217.620 37.490 ;
        RECT 216.610 36.520 216.780 37.320 ;
        RECT 216.985 36.980 217.260 37.120 ;
        RECT 216.980 36.810 217.260 36.980 ;
        RECT 216.265 36.325 216.440 36.360 ;
        RECT 215.510 35.790 215.840 36.190 ;
        RECT 216.265 35.960 216.795 36.325 ;
        RECT 216.985 35.960 217.260 36.810 ;
        RECT 217.430 35.960 217.620 37.320 ;
        RECT 217.790 37.335 217.960 38.000 ;
        RECT 218.130 37.580 218.300 38.340 ;
        RECT 218.535 37.580 219.050 37.990 ;
        RECT 217.790 37.145 218.540 37.335 ;
        RECT 218.710 36.770 219.050 37.580 ;
        RECT 217.820 36.600 219.050 36.770 ;
        RECT 219.220 37.200 219.605 38.170 ;
        RECT 219.775 37.880 220.100 38.340 ;
        RECT 220.620 37.710 220.900 38.170 ;
        RECT 219.775 37.490 220.900 37.710 ;
        RECT 217.800 35.790 218.310 36.325 ;
        RECT 218.530 35.995 218.775 36.600 ;
        RECT 219.220 36.530 219.500 37.200 ;
        RECT 219.775 37.030 220.225 37.490 ;
        RECT 221.090 37.320 221.490 38.170 ;
        RECT 221.890 37.880 222.160 38.340 ;
        RECT 222.330 37.710 222.615 38.170 ;
        RECT 219.670 36.700 220.225 37.030 ;
        RECT 220.395 36.760 221.490 37.320 ;
        RECT 219.775 36.590 220.225 36.700 ;
        RECT 219.220 35.960 219.605 36.530 ;
        RECT 219.775 36.420 220.900 36.590 ;
        RECT 219.775 35.790 220.100 36.250 ;
        RECT 220.620 35.960 220.900 36.420 ;
        RECT 221.090 35.960 221.490 36.760 ;
        RECT 221.660 37.490 222.615 37.710 ;
        RECT 221.660 36.590 221.870 37.490 ;
        RECT 222.040 36.760 222.730 37.320 ;
        RECT 222.900 37.200 223.285 38.170 ;
        RECT 223.455 37.880 223.780 38.340 ;
        RECT 224.300 37.710 224.580 38.170 ;
        RECT 223.455 37.490 224.580 37.710 ;
        RECT 221.660 36.420 222.615 36.590 ;
        RECT 221.890 35.790 222.160 36.250 ;
        RECT 222.330 35.960 222.615 36.420 ;
        RECT 222.900 36.530 223.180 37.200 ;
        RECT 223.455 37.030 223.905 37.490 ;
        RECT 224.770 37.320 225.170 38.170 ;
        RECT 225.570 37.880 225.840 38.340 ;
        RECT 226.010 37.710 226.295 38.170 ;
        RECT 223.350 36.700 223.905 37.030 ;
        RECT 224.075 36.760 225.170 37.320 ;
        RECT 223.455 36.590 223.905 36.700 ;
        RECT 222.900 35.960 223.285 36.530 ;
        RECT 223.455 36.420 224.580 36.590 ;
        RECT 223.455 35.790 223.780 36.250 ;
        RECT 224.300 35.960 224.580 36.420 ;
        RECT 224.770 35.960 225.170 36.760 ;
        RECT 225.340 37.490 226.295 37.710 ;
        RECT 225.340 36.590 225.550 37.490 ;
        RECT 225.720 36.760 226.410 37.320 ;
        RECT 226.580 37.175 226.870 38.340 ;
        RECT 227.040 37.250 228.710 38.340 ;
        RECT 228.885 37.670 229.140 38.170 ;
        RECT 229.310 37.840 229.640 38.340 ;
        RECT 228.885 37.500 229.635 37.670 ;
        RECT 225.340 36.420 226.295 36.590 ;
        RECT 227.040 36.560 227.790 37.080 ;
        RECT 227.960 36.730 228.710 37.250 ;
        RECT 228.885 36.680 229.235 37.330 ;
        RECT 225.570 35.790 225.840 36.250 ;
        RECT 226.010 35.960 226.295 36.420 ;
        RECT 226.580 35.790 226.870 36.515 ;
        RECT 227.040 35.790 228.710 36.560 ;
        RECT 229.405 36.510 229.635 37.500 ;
        RECT 228.885 36.340 229.635 36.510 ;
        RECT 228.885 36.050 229.140 36.340 ;
        RECT 229.310 35.790 229.640 36.170 ;
        RECT 229.810 36.050 229.980 38.170 ;
        RECT 230.150 37.370 230.475 38.155 ;
        RECT 230.645 37.880 230.895 38.340 ;
        RECT 231.065 37.840 231.315 38.170 ;
        RECT 231.530 37.840 232.210 38.170 ;
        RECT 231.065 37.710 231.235 37.840 ;
        RECT 230.840 37.540 231.235 37.710 ;
        RECT 230.210 36.320 230.670 37.370 ;
        RECT 230.840 36.180 231.010 37.540 ;
        RECT 231.405 37.280 231.870 37.670 ;
        RECT 231.180 36.470 231.530 37.090 ;
        RECT 231.700 36.690 231.870 37.280 ;
        RECT 232.040 37.060 232.210 37.840 ;
        RECT 232.380 37.740 232.550 38.080 ;
        RECT 232.785 37.910 233.115 38.340 ;
        RECT 233.285 37.740 233.455 38.080 ;
        RECT 233.750 37.880 234.120 38.340 ;
        RECT 232.380 37.570 233.455 37.740 ;
        RECT 234.290 37.710 234.460 38.170 ;
        RECT 234.695 37.830 235.565 38.170 ;
        RECT 235.735 37.880 235.985 38.340 ;
        RECT 233.900 37.540 234.460 37.710 ;
        RECT 233.900 37.400 234.070 37.540 ;
        RECT 232.570 37.230 234.070 37.400 ;
        RECT 234.765 37.370 235.225 37.660 ;
        RECT 232.040 36.890 233.730 37.060 ;
        RECT 231.700 36.470 232.055 36.690 ;
        RECT 232.225 36.180 232.395 36.890 ;
        RECT 232.600 36.470 233.390 36.720 ;
        RECT 233.560 36.710 233.730 36.890 ;
        RECT 233.900 36.540 234.070 37.230 ;
        RECT 230.340 35.790 230.670 36.150 ;
        RECT 230.840 36.010 231.335 36.180 ;
        RECT 231.540 36.010 232.395 36.180 ;
        RECT 233.270 35.790 233.600 36.250 ;
        RECT 233.810 36.150 234.070 36.540 ;
        RECT 234.260 37.360 235.225 37.370 ;
        RECT 235.395 37.450 235.565 37.830 ;
        RECT 236.155 37.790 236.325 38.080 ;
        RECT 236.505 37.960 236.835 38.340 ;
        RECT 236.155 37.620 236.955 37.790 ;
        RECT 234.260 37.200 234.935 37.360 ;
        RECT 235.395 37.280 236.615 37.450 ;
        RECT 234.260 36.410 234.470 37.200 ;
        RECT 235.395 37.190 235.565 37.280 ;
        RECT 234.640 36.410 234.990 37.030 ;
        RECT 235.160 37.020 235.565 37.190 ;
        RECT 235.160 36.240 235.330 37.020 ;
        RECT 235.500 36.570 235.720 36.850 ;
        RECT 235.900 36.740 236.440 37.110 ;
        RECT 236.785 37.030 236.955 37.620 ;
        RECT 237.175 37.200 237.480 38.340 ;
        RECT 237.650 37.150 237.900 38.030 ;
        RECT 238.070 37.200 238.320 38.340 ;
        RECT 238.540 37.250 239.750 38.340 ;
        RECT 239.925 37.670 240.180 38.170 ;
        RECT 240.350 37.840 240.680 38.340 ;
        RECT 239.925 37.500 240.675 37.670 ;
        RECT 236.785 37.000 237.525 37.030 ;
        RECT 235.500 36.400 236.030 36.570 ;
        RECT 233.810 35.980 234.160 36.150 ;
        RECT 234.380 35.960 235.330 36.240 ;
        RECT 235.500 35.790 235.690 36.230 ;
        RECT 235.860 36.170 236.030 36.400 ;
        RECT 236.200 36.340 236.440 36.740 ;
        RECT 236.610 36.700 237.525 37.000 ;
        RECT 236.610 36.525 236.935 36.700 ;
        RECT 236.610 36.170 236.930 36.525 ;
        RECT 237.695 36.500 237.900 37.150 ;
        RECT 235.860 36.000 236.930 36.170 ;
        RECT 237.175 35.790 237.480 36.250 ;
        RECT 237.650 35.970 237.900 36.500 ;
        RECT 238.070 35.790 238.320 36.545 ;
        RECT 238.540 36.540 239.060 37.080 ;
        RECT 239.230 36.710 239.750 37.250 ;
        RECT 239.925 36.680 240.275 37.330 ;
        RECT 238.540 35.790 239.750 36.540 ;
        RECT 240.445 36.510 240.675 37.500 ;
        RECT 239.925 36.340 240.675 36.510 ;
        RECT 239.925 36.050 240.180 36.340 ;
        RECT 240.350 35.790 240.680 36.170 ;
        RECT 240.850 36.050 241.020 38.170 ;
        RECT 241.190 37.370 241.515 38.155 ;
        RECT 241.685 37.880 241.935 38.340 ;
        RECT 242.105 37.840 242.355 38.170 ;
        RECT 242.570 37.840 243.250 38.170 ;
        RECT 242.105 37.710 242.275 37.840 ;
        RECT 241.880 37.540 242.275 37.710 ;
        RECT 241.250 36.320 241.710 37.370 ;
        RECT 241.880 36.180 242.050 37.540 ;
        RECT 242.445 37.280 242.910 37.670 ;
        RECT 242.220 36.470 242.570 37.090 ;
        RECT 242.740 36.690 242.910 37.280 ;
        RECT 243.080 37.060 243.250 37.840 ;
        RECT 243.420 37.740 243.590 38.080 ;
        RECT 243.825 37.910 244.155 38.340 ;
        RECT 244.325 37.740 244.495 38.080 ;
        RECT 244.790 37.880 245.160 38.340 ;
        RECT 243.420 37.570 244.495 37.740 ;
        RECT 245.330 37.710 245.500 38.170 ;
        RECT 245.735 37.830 246.605 38.170 ;
        RECT 246.775 37.880 247.025 38.340 ;
        RECT 244.940 37.540 245.500 37.710 ;
        RECT 244.940 37.400 245.110 37.540 ;
        RECT 243.610 37.230 245.110 37.400 ;
        RECT 245.805 37.370 246.265 37.660 ;
        RECT 243.080 36.890 244.770 37.060 ;
        RECT 242.740 36.470 243.095 36.690 ;
        RECT 243.265 36.180 243.435 36.890 ;
        RECT 243.640 36.470 244.430 36.720 ;
        RECT 244.600 36.710 244.770 36.890 ;
        RECT 244.940 36.540 245.110 37.230 ;
        RECT 241.380 35.790 241.710 36.150 ;
        RECT 241.880 36.010 242.375 36.180 ;
        RECT 242.580 36.010 243.435 36.180 ;
        RECT 244.310 35.790 244.640 36.250 ;
        RECT 244.850 36.150 245.110 36.540 ;
        RECT 245.300 37.360 246.265 37.370 ;
        RECT 246.435 37.450 246.605 37.830 ;
        RECT 247.195 37.790 247.365 38.080 ;
        RECT 247.545 37.960 247.875 38.340 ;
        RECT 247.195 37.620 247.995 37.790 ;
        RECT 245.300 37.200 245.975 37.360 ;
        RECT 246.435 37.280 247.655 37.450 ;
        RECT 245.300 36.410 245.510 37.200 ;
        RECT 246.435 37.190 246.605 37.280 ;
        RECT 245.680 36.410 246.030 37.030 ;
        RECT 246.200 37.020 246.605 37.190 ;
        RECT 246.200 36.240 246.370 37.020 ;
        RECT 246.540 36.570 246.760 36.850 ;
        RECT 246.940 36.740 247.480 37.110 ;
        RECT 247.825 37.030 247.995 37.620 ;
        RECT 248.215 37.200 248.520 38.340 ;
        RECT 248.690 37.150 248.945 38.030 ;
        RECT 249.120 37.250 251.710 38.340 ;
        RECT 247.825 37.000 248.565 37.030 ;
        RECT 246.540 36.400 247.070 36.570 ;
        RECT 244.850 35.980 245.200 36.150 ;
        RECT 245.420 35.960 246.370 36.240 ;
        RECT 246.540 35.790 246.730 36.230 ;
        RECT 246.900 36.170 247.070 36.400 ;
        RECT 247.240 36.340 247.480 36.740 ;
        RECT 247.650 36.700 248.565 37.000 ;
        RECT 247.650 36.525 247.975 36.700 ;
        RECT 247.650 36.170 247.970 36.525 ;
        RECT 248.735 36.500 248.945 37.150 ;
        RECT 246.900 36.000 247.970 36.170 ;
        RECT 248.215 35.790 248.520 36.250 ;
        RECT 248.690 35.970 248.945 36.500 ;
        RECT 249.120 36.560 250.330 37.080 ;
        RECT 250.500 36.730 251.710 37.250 ;
        RECT 252.340 37.175 252.630 38.340 ;
        RECT 252.800 37.250 254.010 38.340 ;
        RECT 254.185 37.670 254.440 38.170 ;
        RECT 254.610 37.840 254.940 38.340 ;
        RECT 254.185 37.500 254.935 37.670 ;
        RECT 249.120 35.790 251.710 36.560 ;
        RECT 252.800 36.540 253.320 37.080 ;
        RECT 253.490 36.710 254.010 37.250 ;
        RECT 254.185 36.680 254.535 37.330 ;
        RECT 252.340 35.790 252.630 36.515 ;
        RECT 252.800 35.790 254.010 36.540 ;
        RECT 254.705 36.510 254.935 37.500 ;
        RECT 254.185 36.340 254.935 36.510 ;
        RECT 254.185 36.050 254.440 36.340 ;
        RECT 254.610 35.790 254.940 36.170 ;
        RECT 255.110 36.050 255.280 38.170 ;
        RECT 255.450 37.370 255.775 38.155 ;
        RECT 255.945 37.880 256.195 38.340 ;
        RECT 256.365 37.840 256.615 38.170 ;
        RECT 256.830 37.840 257.510 38.170 ;
        RECT 256.365 37.710 256.535 37.840 ;
        RECT 256.140 37.540 256.535 37.710 ;
        RECT 255.510 36.320 255.970 37.370 ;
        RECT 256.140 36.180 256.310 37.540 ;
        RECT 256.705 37.280 257.170 37.670 ;
        RECT 256.480 36.470 256.830 37.090 ;
        RECT 257.000 36.690 257.170 37.280 ;
        RECT 257.340 37.060 257.510 37.840 ;
        RECT 257.680 37.740 257.850 38.080 ;
        RECT 258.085 37.910 258.415 38.340 ;
        RECT 258.585 37.740 258.755 38.080 ;
        RECT 259.050 37.880 259.420 38.340 ;
        RECT 257.680 37.570 258.755 37.740 ;
        RECT 259.590 37.710 259.760 38.170 ;
        RECT 259.995 37.830 260.865 38.170 ;
        RECT 261.035 37.880 261.285 38.340 ;
        RECT 259.200 37.540 259.760 37.710 ;
        RECT 259.200 37.400 259.370 37.540 ;
        RECT 257.870 37.230 259.370 37.400 ;
        RECT 260.065 37.370 260.525 37.660 ;
        RECT 257.340 36.890 259.030 37.060 ;
        RECT 257.000 36.470 257.355 36.690 ;
        RECT 257.525 36.180 257.695 36.890 ;
        RECT 257.900 36.470 258.690 36.720 ;
        RECT 258.860 36.710 259.030 36.890 ;
        RECT 259.200 36.540 259.370 37.230 ;
        RECT 255.640 35.790 255.970 36.150 ;
        RECT 256.140 36.010 256.635 36.180 ;
        RECT 256.840 36.010 257.695 36.180 ;
        RECT 258.570 35.790 258.900 36.250 ;
        RECT 259.110 36.150 259.370 36.540 ;
        RECT 259.560 37.360 260.525 37.370 ;
        RECT 260.695 37.450 260.865 37.830 ;
        RECT 261.455 37.790 261.625 38.080 ;
        RECT 261.805 37.960 262.135 38.340 ;
        RECT 261.455 37.620 262.255 37.790 ;
        RECT 259.560 37.200 260.235 37.360 ;
        RECT 260.695 37.280 261.915 37.450 ;
        RECT 259.560 36.410 259.770 37.200 ;
        RECT 260.695 37.190 260.865 37.280 ;
        RECT 259.940 36.410 260.290 37.030 ;
        RECT 260.460 37.020 260.865 37.190 ;
        RECT 260.460 36.240 260.630 37.020 ;
        RECT 260.800 36.570 261.020 36.850 ;
        RECT 261.200 36.740 261.740 37.110 ;
        RECT 262.085 37.030 262.255 37.620 ;
        RECT 262.475 37.200 262.780 38.340 ;
        RECT 262.950 37.150 263.205 38.030 ;
        RECT 262.085 37.000 262.825 37.030 ;
        RECT 260.800 36.400 261.330 36.570 ;
        RECT 259.110 35.980 259.460 36.150 ;
        RECT 259.680 35.960 260.630 36.240 ;
        RECT 260.800 35.790 260.990 36.230 ;
        RECT 261.160 36.170 261.330 36.400 ;
        RECT 261.500 36.340 261.740 36.740 ;
        RECT 261.910 36.700 262.825 37.000 ;
        RECT 261.910 36.525 262.235 36.700 ;
        RECT 261.910 36.170 262.230 36.525 ;
        RECT 262.995 36.500 263.205 37.150 ;
        RECT 261.160 36.000 262.230 36.170 ;
        RECT 262.475 35.790 262.780 36.250 ;
        RECT 262.950 35.970 263.205 36.500 ;
        RECT 263.415 37.550 263.950 38.170 ;
        RECT 263.415 36.530 263.730 37.550 ;
        RECT 264.120 37.540 264.450 38.340 ;
        RECT 265.680 37.620 266.140 38.170 ;
        RECT 266.330 37.620 266.660 38.340 ;
        RECT 264.935 37.370 265.325 37.545 ;
        RECT 263.900 37.200 265.325 37.370 ;
        RECT 263.900 36.700 264.070 37.200 ;
        RECT 263.415 35.960 264.030 36.530 ;
        RECT 264.320 36.470 264.585 37.030 ;
        RECT 264.755 36.300 264.925 37.200 ;
        RECT 265.095 36.470 265.450 37.030 ;
        RECT 264.200 35.790 264.415 36.300 ;
        RECT 264.645 35.970 264.925 36.300 ;
        RECT 265.105 35.790 265.345 36.300 ;
        RECT 265.680 36.250 265.930 37.620 ;
        RECT 266.860 37.450 267.160 38.000 ;
        RECT 267.330 37.670 267.610 38.340 ;
        RECT 268.905 37.670 269.160 38.170 ;
        RECT 269.330 37.840 269.660 38.340 ;
        RECT 268.905 37.500 269.655 37.670 ;
        RECT 266.220 37.280 267.160 37.450 ;
        RECT 266.220 37.030 266.390 37.280 ;
        RECT 267.530 37.030 267.795 37.390 ;
        RECT 266.100 36.700 266.390 37.030 ;
        RECT 266.560 36.780 266.900 37.030 ;
        RECT 267.120 36.780 267.795 37.030 ;
        RECT 266.220 36.610 266.390 36.700 ;
        RECT 268.905 36.680 269.255 37.330 ;
        RECT 266.220 36.420 267.610 36.610 ;
        RECT 269.425 36.510 269.655 37.500 ;
        RECT 265.680 35.960 266.240 36.250 ;
        RECT 266.410 35.790 266.660 36.250 ;
        RECT 267.280 36.060 267.610 36.420 ;
        RECT 268.905 36.340 269.655 36.510 ;
        RECT 268.905 36.050 269.160 36.340 ;
        RECT 269.330 35.790 269.660 36.170 ;
        RECT 269.830 36.050 270.000 38.170 ;
        RECT 270.170 37.370 270.495 38.155 ;
        RECT 270.665 37.880 270.915 38.340 ;
        RECT 271.085 37.840 271.335 38.170 ;
        RECT 271.550 37.840 272.230 38.170 ;
        RECT 271.085 37.710 271.255 37.840 ;
        RECT 270.860 37.540 271.255 37.710 ;
        RECT 270.230 36.320 270.690 37.370 ;
        RECT 270.860 36.180 271.030 37.540 ;
        RECT 271.425 37.280 271.890 37.670 ;
        RECT 271.200 36.470 271.550 37.090 ;
        RECT 271.720 36.690 271.890 37.280 ;
        RECT 272.060 37.060 272.230 37.840 ;
        RECT 272.400 37.740 272.570 38.080 ;
        RECT 272.805 37.910 273.135 38.340 ;
        RECT 273.305 37.740 273.475 38.080 ;
        RECT 273.770 37.880 274.140 38.340 ;
        RECT 272.400 37.570 273.475 37.740 ;
        RECT 274.310 37.710 274.480 38.170 ;
        RECT 274.715 37.830 275.585 38.170 ;
        RECT 275.755 37.880 276.005 38.340 ;
        RECT 273.920 37.540 274.480 37.710 ;
        RECT 273.920 37.400 274.090 37.540 ;
        RECT 272.590 37.230 274.090 37.400 ;
        RECT 274.785 37.370 275.245 37.660 ;
        RECT 272.060 36.890 273.750 37.060 ;
        RECT 271.720 36.470 272.075 36.690 ;
        RECT 272.245 36.180 272.415 36.890 ;
        RECT 272.620 36.470 273.410 36.720 ;
        RECT 273.580 36.710 273.750 36.890 ;
        RECT 273.920 36.540 274.090 37.230 ;
        RECT 270.360 35.790 270.690 36.150 ;
        RECT 270.860 36.010 271.355 36.180 ;
        RECT 271.560 36.010 272.415 36.180 ;
        RECT 273.290 35.790 273.620 36.250 ;
        RECT 273.830 36.150 274.090 36.540 ;
        RECT 274.280 37.360 275.245 37.370 ;
        RECT 275.415 37.450 275.585 37.830 ;
        RECT 276.175 37.790 276.345 38.080 ;
        RECT 276.525 37.960 276.855 38.340 ;
        RECT 276.175 37.620 276.975 37.790 ;
        RECT 274.280 37.200 274.955 37.360 ;
        RECT 275.415 37.280 276.635 37.450 ;
        RECT 274.280 36.410 274.490 37.200 ;
        RECT 275.415 37.190 275.585 37.280 ;
        RECT 274.660 36.410 275.010 37.030 ;
        RECT 275.180 37.020 275.585 37.190 ;
        RECT 275.180 36.240 275.350 37.020 ;
        RECT 275.520 36.570 275.740 36.850 ;
        RECT 275.920 36.740 276.460 37.110 ;
        RECT 276.805 37.030 276.975 37.620 ;
        RECT 277.195 37.200 277.500 38.340 ;
        RECT 277.670 37.150 277.925 38.030 ;
        RECT 278.100 37.175 278.390 38.340 ;
        RECT 278.560 37.830 278.820 38.340 ;
        RECT 276.805 37.000 277.545 37.030 ;
        RECT 275.520 36.400 276.050 36.570 ;
        RECT 273.830 35.980 274.180 36.150 ;
        RECT 274.400 35.960 275.350 36.240 ;
        RECT 275.520 35.790 275.710 36.230 ;
        RECT 275.880 36.170 276.050 36.400 ;
        RECT 276.220 36.340 276.460 36.740 ;
        RECT 276.630 36.700 277.545 37.000 ;
        RECT 276.630 36.525 276.955 36.700 ;
        RECT 276.630 36.170 276.950 36.525 ;
        RECT 277.715 36.500 277.925 37.150 ;
        RECT 278.560 36.780 278.900 37.660 ;
        RECT 279.070 36.950 279.240 38.170 ;
        RECT 279.480 37.835 280.095 38.340 ;
        RECT 279.480 37.300 279.730 37.665 ;
        RECT 279.900 37.660 280.095 37.835 ;
        RECT 280.265 37.830 280.740 38.170 ;
        RECT 280.910 37.795 281.125 38.340 ;
        RECT 279.900 37.470 280.230 37.660 ;
        RECT 280.450 37.300 281.165 37.595 ;
        RECT 281.335 37.470 281.610 38.170 ;
        RECT 281.780 37.905 287.125 38.340 ;
        RECT 287.300 37.905 292.645 38.340 ;
        RECT 292.820 37.905 298.165 38.340 ;
        RECT 298.340 37.905 303.685 38.340 ;
        RECT 279.480 37.130 281.270 37.300 ;
        RECT 279.070 36.700 279.865 36.950 ;
        RECT 279.070 36.610 279.320 36.700 ;
        RECT 275.880 36.000 276.950 36.170 ;
        RECT 277.195 35.790 277.500 36.250 ;
        RECT 277.670 35.970 277.925 36.500 ;
        RECT 278.100 35.790 278.390 36.515 ;
        RECT 278.560 35.790 278.820 36.610 ;
        RECT 278.990 36.190 279.320 36.610 ;
        RECT 280.035 36.275 280.290 37.130 ;
        RECT 279.500 36.010 280.290 36.275 ;
        RECT 280.460 36.430 280.870 36.950 ;
        RECT 281.040 36.700 281.270 37.130 ;
        RECT 281.440 36.440 281.610 37.470 ;
        RECT 280.460 36.010 280.660 36.430 ;
        RECT 280.850 35.790 281.180 36.250 ;
        RECT 281.350 35.960 281.610 36.440 ;
        RECT 283.365 36.335 283.705 37.165 ;
        RECT 285.185 36.655 285.535 37.905 ;
        RECT 288.885 36.335 289.225 37.165 ;
        RECT 290.705 36.655 291.055 37.905 ;
        RECT 294.405 36.335 294.745 37.165 ;
        RECT 296.225 36.655 296.575 37.905 ;
        RECT 299.925 36.335 300.265 37.165 ;
        RECT 301.745 36.655 302.095 37.905 ;
        RECT 303.860 37.175 304.150 38.340 ;
        RECT 304.320 37.250 307.830 38.340 ;
        RECT 308.005 37.915 308.340 38.340 ;
        RECT 308.510 37.735 308.695 38.140 ;
        RECT 304.320 36.560 305.970 37.080 ;
        RECT 306.140 36.730 307.830 37.250 ;
        RECT 308.030 37.560 308.695 37.735 ;
        RECT 308.900 37.560 309.230 38.340 ;
        RECT 281.780 35.790 287.125 36.335 ;
        RECT 287.300 35.790 292.645 36.335 ;
        RECT 292.820 35.790 298.165 36.335 ;
        RECT 298.340 35.790 303.685 36.335 ;
        RECT 303.860 35.790 304.150 36.515 ;
        RECT 304.320 35.790 307.830 36.560 ;
        RECT 308.030 36.530 308.370 37.560 ;
        RECT 309.400 37.370 309.670 38.140 ;
        RECT 308.540 37.200 309.670 37.370 ;
        RECT 308.540 36.700 308.790 37.200 ;
        RECT 308.030 36.360 308.715 36.530 ;
        RECT 308.970 36.450 309.330 37.030 ;
        RECT 308.005 35.790 308.340 36.190 ;
        RECT 308.510 35.960 308.715 36.360 ;
        RECT 309.500 36.290 309.670 37.200 ;
        RECT 309.840 37.250 311.050 38.340 ;
        RECT 309.840 36.710 310.360 37.250 ;
        RECT 310.530 36.540 311.050 37.080 ;
        RECT 308.925 35.790 309.200 36.270 ;
        RECT 309.410 35.960 309.670 36.290 ;
        RECT 309.840 35.790 311.050 36.540 ;
        RECT 162.095 35.620 311.135 35.790 ;
        RECT 162.180 34.870 163.390 35.620 ;
        RECT 162.180 34.330 162.700 34.870 ;
        RECT 163.560 34.850 165.230 35.620 ;
        RECT 165.865 35.070 166.120 35.360 ;
        RECT 166.290 35.240 166.620 35.620 ;
        RECT 165.865 34.900 166.615 35.070 ;
        RECT 162.870 34.160 163.390 34.700 ;
        RECT 163.560 34.330 164.310 34.850 ;
        RECT 164.480 34.160 165.230 34.680 ;
        RECT 162.180 33.070 163.390 34.160 ;
        RECT 163.560 33.070 165.230 34.160 ;
        RECT 165.865 34.080 166.215 34.730 ;
        RECT 166.385 33.910 166.615 34.900 ;
        RECT 165.865 33.740 166.615 33.910 ;
        RECT 165.865 33.240 166.120 33.740 ;
        RECT 166.290 33.070 166.620 33.570 ;
        RECT 166.790 33.240 166.960 35.360 ;
        RECT 167.320 35.260 167.650 35.620 ;
        RECT 167.820 35.230 168.315 35.400 ;
        RECT 168.520 35.230 169.375 35.400 ;
        RECT 167.190 34.040 167.650 35.090 ;
        RECT 167.130 33.255 167.455 34.040 ;
        RECT 167.820 33.870 167.990 35.230 ;
        RECT 168.160 34.320 168.510 34.940 ;
        RECT 168.680 34.720 169.035 34.940 ;
        RECT 168.680 34.130 168.850 34.720 ;
        RECT 169.205 34.520 169.375 35.230 ;
        RECT 170.250 35.160 170.580 35.620 ;
        RECT 170.790 35.260 171.140 35.430 ;
        RECT 169.580 34.690 170.370 34.940 ;
        RECT 170.790 34.870 171.050 35.260 ;
        RECT 171.360 35.170 172.310 35.450 ;
        RECT 172.480 35.180 172.670 35.620 ;
        RECT 172.840 35.240 173.910 35.410 ;
        RECT 170.540 34.520 170.710 34.700 ;
        RECT 167.820 33.700 168.215 33.870 ;
        RECT 168.385 33.740 168.850 34.130 ;
        RECT 169.020 34.350 170.710 34.520 ;
        RECT 168.045 33.570 168.215 33.700 ;
        RECT 169.020 33.570 169.190 34.350 ;
        RECT 170.880 34.180 171.050 34.870 ;
        RECT 169.550 34.010 171.050 34.180 ;
        RECT 171.240 34.210 171.450 35.000 ;
        RECT 171.620 34.380 171.970 35.000 ;
        RECT 172.140 34.390 172.310 35.170 ;
        RECT 172.840 35.010 173.010 35.240 ;
        RECT 172.480 34.840 173.010 35.010 ;
        RECT 172.480 34.560 172.700 34.840 ;
        RECT 173.180 34.670 173.420 35.070 ;
        RECT 172.140 34.220 172.545 34.390 ;
        RECT 172.880 34.300 173.420 34.670 ;
        RECT 173.590 34.885 173.910 35.240 ;
        RECT 174.155 35.160 174.460 35.620 ;
        RECT 174.630 34.910 174.885 35.440 ;
        RECT 173.590 34.710 173.915 34.885 ;
        RECT 173.590 34.410 174.505 34.710 ;
        RECT 173.765 34.380 174.505 34.410 ;
        RECT 171.240 34.050 171.915 34.210 ;
        RECT 172.375 34.130 172.545 34.220 ;
        RECT 171.240 34.040 172.205 34.050 ;
        RECT 170.880 33.870 171.050 34.010 ;
        RECT 167.625 33.070 167.875 33.530 ;
        RECT 168.045 33.240 168.295 33.570 ;
        RECT 168.510 33.240 169.190 33.570 ;
        RECT 169.360 33.670 170.435 33.840 ;
        RECT 170.880 33.700 171.440 33.870 ;
        RECT 171.745 33.750 172.205 34.040 ;
        RECT 172.375 33.960 173.595 34.130 ;
        RECT 169.360 33.330 169.530 33.670 ;
        RECT 169.765 33.070 170.095 33.500 ;
        RECT 170.265 33.330 170.435 33.670 ;
        RECT 170.730 33.070 171.100 33.530 ;
        RECT 171.270 33.240 171.440 33.700 ;
        RECT 172.375 33.580 172.545 33.960 ;
        RECT 173.765 33.790 173.935 34.380 ;
        RECT 174.675 34.260 174.885 34.910 ;
        RECT 171.675 33.240 172.545 33.580 ;
        RECT 173.135 33.620 173.935 33.790 ;
        RECT 172.715 33.070 172.965 33.530 ;
        RECT 173.135 33.330 173.305 33.620 ;
        RECT 173.485 33.070 173.815 33.450 ;
        RECT 174.155 33.070 174.460 34.210 ;
        RECT 174.630 33.380 174.885 34.260 ;
        RECT 175.060 34.880 175.445 35.450 ;
        RECT 175.615 35.160 175.940 35.620 ;
        RECT 176.460 34.990 176.740 35.450 ;
        RECT 175.060 34.210 175.340 34.880 ;
        RECT 175.615 34.820 176.740 34.990 ;
        RECT 175.615 34.710 176.065 34.820 ;
        RECT 175.510 34.380 176.065 34.710 ;
        RECT 176.930 34.650 177.330 35.450 ;
        RECT 177.730 35.160 178.000 35.620 ;
        RECT 178.170 34.990 178.455 35.450 ;
        RECT 175.060 33.240 175.445 34.210 ;
        RECT 175.615 33.920 176.065 34.380 ;
        RECT 176.235 34.090 177.330 34.650 ;
        RECT 175.615 33.700 176.740 33.920 ;
        RECT 175.615 33.070 175.940 33.530 ;
        RECT 176.460 33.240 176.740 33.700 ;
        RECT 176.930 33.240 177.330 34.090 ;
        RECT 177.500 34.820 178.455 34.990 ;
        RECT 178.745 34.910 179.000 35.440 ;
        RECT 179.170 35.160 179.475 35.620 ;
        RECT 179.720 35.240 180.790 35.410 ;
        RECT 177.500 33.920 177.710 34.820 ;
        RECT 177.880 34.090 178.570 34.650 ;
        RECT 178.745 34.260 178.955 34.910 ;
        RECT 179.720 34.885 180.040 35.240 ;
        RECT 179.715 34.710 180.040 34.885 ;
        RECT 179.125 34.410 180.040 34.710 ;
        RECT 180.210 34.670 180.450 35.070 ;
        RECT 180.620 35.010 180.790 35.240 ;
        RECT 180.960 35.180 181.150 35.620 ;
        RECT 181.320 35.170 182.270 35.450 ;
        RECT 182.490 35.260 182.840 35.430 ;
        RECT 180.620 34.840 181.150 35.010 ;
        RECT 179.125 34.380 179.865 34.410 ;
        RECT 177.500 33.700 178.455 33.920 ;
        RECT 177.730 33.070 178.000 33.530 ;
        RECT 178.170 33.240 178.455 33.700 ;
        RECT 178.745 33.380 179.000 34.260 ;
        RECT 179.170 33.070 179.475 34.210 ;
        RECT 179.695 33.790 179.865 34.380 ;
        RECT 180.210 34.300 180.750 34.670 ;
        RECT 180.930 34.560 181.150 34.840 ;
        RECT 181.320 34.390 181.490 35.170 ;
        RECT 181.085 34.220 181.490 34.390 ;
        RECT 181.660 34.380 182.010 35.000 ;
        RECT 181.085 34.130 181.255 34.220 ;
        RECT 182.180 34.210 182.390 35.000 ;
        RECT 180.035 33.960 181.255 34.130 ;
        RECT 181.715 34.050 182.390 34.210 ;
        RECT 179.695 33.620 180.495 33.790 ;
        RECT 179.815 33.070 180.145 33.450 ;
        RECT 180.325 33.330 180.495 33.620 ;
        RECT 181.085 33.580 181.255 33.960 ;
        RECT 181.425 34.040 182.390 34.050 ;
        RECT 182.580 34.870 182.840 35.260 ;
        RECT 183.050 35.160 183.380 35.620 ;
        RECT 184.255 35.230 185.110 35.400 ;
        RECT 185.315 35.230 185.810 35.400 ;
        RECT 185.980 35.260 186.310 35.620 ;
        RECT 182.580 34.180 182.750 34.870 ;
        RECT 182.920 34.520 183.090 34.700 ;
        RECT 183.260 34.690 184.050 34.940 ;
        RECT 184.255 34.520 184.425 35.230 ;
        RECT 184.595 34.720 184.950 34.940 ;
        RECT 182.920 34.350 184.610 34.520 ;
        RECT 181.425 33.750 181.885 34.040 ;
        RECT 182.580 34.010 184.080 34.180 ;
        RECT 182.580 33.870 182.750 34.010 ;
        RECT 182.190 33.700 182.750 33.870 ;
        RECT 180.665 33.070 180.915 33.530 ;
        RECT 181.085 33.240 181.955 33.580 ;
        RECT 182.190 33.240 182.360 33.700 ;
        RECT 183.195 33.670 184.270 33.840 ;
        RECT 182.530 33.070 182.900 33.530 ;
        RECT 183.195 33.330 183.365 33.670 ;
        RECT 183.535 33.070 183.865 33.500 ;
        RECT 184.100 33.330 184.270 33.670 ;
        RECT 184.440 33.570 184.610 34.350 ;
        RECT 184.780 34.130 184.950 34.720 ;
        RECT 185.120 34.320 185.470 34.940 ;
        RECT 184.780 33.740 185.245 34.130 ;
        RECT 185.640 33.870 185.810 35.230 ;
        RECT 185.980 34.040 186.440 35.090 ;
        RECT 185.415 33.700 185.810 33.870 ;
        RECT 185.415 33.570 185.585 33.700 ;
        RECT 184.440 33.240 185.120 33.570 ;
        RECT 185.335 33.240 185.585 33.570 ;
        RECT 185.755 33.070 186.005 33.530 ;
        RECT 186.175 33.255 186.500 34.040 ;
        RECT 186.670 33.240 186.840 35.360 ;
        RECT 187.010 35.240 187.340 35.620 ;
        RECT 187.510 35.070 187.765 35.360 ;
        RECT 187.015 34.900 187.765 35.070 ;
        RECT 187.015 33.910 187.245 34.900 ;
        RECT 187.940 34.895 188.230 35.620 ;
        RECT 188.405 35.070 188.660 35.360 ;
        RECT 188.830 35.240 189.160 35.620 ;
        RECT 188.405 34.900 189.155 35.070 ;
        RECT 187.415 34.080 187.765 34.730 ;
        RECT 187.015 33.740 187.765 33.910 ;
        RECT 187.010 33.070 187.340 33.570 ;
        RECT 187.510 33.240 187.765 33.740 ;
        RECT 187.940 33.070 188.230 34.235 ;
        RECT 188.405 34.080 188.755 34.730 ;
        RECT 188.925 33.910 189.155 34.900 ;
        RECT 188.405 33.740 189.155 33.910 ;
        RECT 188.405 33.240 188.660 33.740 ;
        RECT 188.830 33.070 189.160 33.570 ;
        RECT 189.330 33.240 189.500 35.360 ;
        RECT 189.860 35.260 190.190 35.620 ;
        RECT 190.360 35.230 190.855 35.400 ;
        RECT 191.060 35.230 191.915 35.400 ;
        RECT 189.730 34.040 190.190 35.090 ;
        RECT 189.670 33.255 189.995 34.040 ;
        RECT 190.360 33.870 190.530 35.230 ;
        RECT 190.700 34.320 191.050 34.940 ;
        RECT 191.220 34.720 191.575 34.940 ;
        RECT 191.220 34.130 191.390 34.720 ;
        RECT 191.745 34.520 191.915 35.230 ;
        RECT 192.790 35.160 193.120 35.620 ;
        RECT 193.330 35.260 193.680 35.430 ;
        RECT 192.120 34.690 192.910 34.940 ;
        RECT 193.330 34.870 193.590 35.260 ;
        RECT 193.900 35.170 194.850 35.450 ;
        RECT 195.020 35.180 195.210 35.620 ;
        RECT 195.380 35.240 196.450 35.410 ;
        RECT 193.080 34.520 193.250 34.700 ;
        RECT 190.360 33.700 190.755 33.870 ;
        RECT 190.925 33.740 191.390 34.130 ;
        RECT 191.560 34.350 193.250 34.520 ;
        RECT 190.585 33.570 190.755 33.700 ;
        RECT 191.560 33.570 191.730 34.350 ;
        RECT 193.420 34.180 193.590 34.870 ;
        RECT 192.090 34.010 193.590 34.180 ;
        RECT 193.780 34.210 193.990 35.000 ;
        RECT 194.160 34.380 194.510 35.000 ;
        RECT 194.680 34.390 194.850 35.170 ;
        RECT 195.380 35.010 195.550 35.240 ;
        RECT 195.020 34.840 195.550 35.010 ;
        RECT 195.020 34.560 195.240 34.840 ;
        RECT 195.720 34.670 195.960 35.070 ;
        RECT 194.680 34.220 195.085 34.390 ;
        RECT 195.420 34.300 195.960 34.670 ;
        RECT 196.130 34.885 196.450 35.240 ;
        RECT 196.695 35.160 197.000 35.620 ;
        RECT 197.170 34.910 197.425 35.440 ;
        RECT 196.130 34.710 196.455 34.885 ;
        RECT 196.130 34.410 197.045 34.710 ;
        RECT 196.305 34.380 197.045 34.410 ;
        RECT 193.780 34.050 194.455 34.210 ;
        RECT 194.915 34.130 195.085 34.220 ;
        RECT 193.780 34.040 194.745 34.050 ;
        RECT 193.420 33.870 193.590 34.010 ;
        RECT 190.165 33.070 190.415 33.530 ;
        RECT 190.585 33.240 190.835 33.570 ;
        RECT 191.050 33.240 191.730 33.570 ;
        RECT 191.900 33.670 192.975 33.840 ;
        RECT 193.420 33.700 193.980 33.870 ;
        RECT 194.285 33.750 194.745 34.040 ;
        RECT 194.915 33.960 196.135 34.130 ;
        RECT 191.900 33.330 192.070 33.670 ;
        RECT 192.305 33.070 192.635 33.500 ;
        RECT 192.805 33.330 192.975 33.670 ;
        RECT 193.270 33.070 193.640 33.530 ;
        RECT 193.810 33.240 193.980 33.700 ;
        RECT 194.915 33.580 195.085 33.960 ;
        RECT 196.305 33.790 196.475 34.380 ;
        RECT 197.215 34.260 197.425 34.910 ;
        RECT 194.215 33.240 195.085 33.580 ;
        RECT 195.675 33.620 196.475 33.790 ;
        RECT 195.255 33.070 195.505 33.530 ;
        RECT 195.675 33.330 195.845 33.620 ;
        RECT 196.025 33.070 196.355 33.450 ;
        RECT 196.695 33.070 197.000 34.210 ;
        RECT 197.170 33.380 197.425 34.260 ;
        RECT 197.600 34.880 197.985 35.450 ;
        RECT 198.155 35.160 198.480 35.620 ;
        RECT 199.000 34.990 199.280 35.450 ;
        RECT 197.600 34.210 197.880 34.880 ;
        RECT 198.155 34.820 199.280 34.990 ;
        RECT 198.155 34.710 198.605 34.820 ;
        RECT 198.050 34.380 198.605 34.710 ;
        RECT 199.470 34.650 199.870 35.450 ;
        RECT 200.270 35.160 200.540 35.620 ;
        RECT 200.710 34.990 200.995 35.450 ;
        RECT 197.600 33.240 197.985 34.210 ;
        RECT 198.155 33.920 198.605 34.380 ;
        RECT 198.775 34.090 199.870 34.650 ;
        RECT 198.155 33.700 199.280 33.920 ;
        RECT 198.155 33.070 198.480 33.530 ;
        RECT 199.000 33.240 199.280 33.700 ;
        RECT 199.470 33.240 199.870 34.090 ;
        RECT 200.040 34.820 200.995 34.990 ;
        RECT 201.285 35.070 201.540 35.360 ;
        RECT 201.710 35.240 202.040 35.620 ;
        RECT 201.285 34.900 202.035 35.070 ;
        RECT 200.040 33.920 200.250 34.820 ;
        RECT 200.420 34.090 201.110 34.650 ;
        RECT 201.285 34.080 201.635 34.730 ;
        RECT 200.040 33.700 200.995 33.920 ;
        RECT 201.805 33.910 202.035 34.900 ;
        RECT 200.270 33.070 200.540 33.530 ;
        RECT 200.710 33.240 200.995 33.700 ;
        RECT 201.285 33.740 202.035 33.910 ;
        RECT 201.285 33.240 201.540 33.740 ;
        RECT 201.710 33.070 202.040 33.570 ;
        RECT 202.210 33.240 202.380 35.360 ;
        RECT 202.740 35.260 203.070 35.620 ;
        RECT 203.240 35.230 203.735 35.400 ;
        RECT 203.940 35.230 204.795 35.400 ;
        RECT 202.610 34.040 203.070 35.090 ;
        RECT 202.550 33.255 202.875 34.040 ;
        RECT 203.240 33.870 203.410 35.230 ;
        RECT 203.580 34.320 203.930 34.940 ;
        RECT 204.100 34.720 204.455 34.940 ;
        RECT 204.100 34.130 204.270 34.720 ;
        RECT 204.625 34.520 204.795 35.230 ;
        RECT 205.670 35.160 206.000 35.620 ;
        RECT 206.210 35.260 206.560 35.430 ;
        RECT 205.000 34.690 205.790 34.940 ;
        RECT 206.210 34.870 206.470 35.260 ;
        RECT 206.780 35.170 207.730 35.450 ;
        RECT 207.900 35.180 208.090 35.620 ;
        RECT 208.260 35.240 209.330 35.410 ;
        RECT 205.960 34.520 206.130 34.700 ;
        RECT 203.240 33.700 203.635 33.870 ;
        RECT 203.805 33.740 204.270 34.130 ;
        RECT 204.440 34.350 206.130 34.520 ;
        RECT 203.465 33.570 203.635 33.700 ;
        RECT 204.440 33.570 204.610 34.350 ;
        RECT 206.300 34.180 206.470 34.870 ;
        RECT 204.970 34.010 206.470 34.180 ;
        RECT 206.660 34.210 206.870 35.000 ;
        RECT 207.040 34.380 207.390 35.000 ;
        RECT 207.560 34.390 207.730 35.170 ;
        RECT 208.260 35.010 208.430 35.240 ;
        RECT 207.900 34.840 208.430 35.010 ;
        RECT 207.900 34.560 208.120 34.840 ;
        RECT 208.600 34.670 208.840 35.070 ;
        RECT 207.560 34.220 207.965 34.390 ;
        RECT 208.300 34.300 208.840 34.670 ;
        RECT 209.010 34.885 209.330 35.240 ;
        RECT 209.575 35.160 209.880 35.620 ;
        RECT 210.050 34.910 210.305 35.440 ;
        RECT 210.540 35.140 210.820 35.620 ;
        RECT 210.990 34.970 211.250 35.360 ;
        RECT 211.425 35.140 211.680 35.620 ;
        RECT 211.850 34.970 212.145 35.360 ;
        RECT 212.325 35.140 212.600 35.620 ;
        RECT 212.770 35.120 213.070 35.450 ;
        RECT 209.010 34.710 209.335 34.885 ;
        RECT 209.010 34.410 209.925 34.710 ;
        RECT 209.185 34.380 209.925 34.410 ;
        RECT 206.660 34.050 207.335 34.210 ;
        RECT 207.795 34.130 207.965 34.220 ;
        RECT 206.660 34.040 207.625 34.050 ;
        RECT 206.300 33.870 206.470 34.010 ;
        RECT 203.045 33.070 203.295 33.530 ;
        RECT 203.465 33.240 203.715 33.570 ;
        RECT 203.930 33.240 204.610 33.570 ;
        RECT 204.780 33.670 205.855 33.840 ;
        RECT 206.300 33.700 206.860 33.870 ;
        RECT 207.165 33.750 207.625 34.040 ;
        RECT 207.795 33.960 209.015 34.130 ;
        RECT 204.780 33.330 204.950 33.670 ;
        RECT 205.185 33.070 205.515 33.500 ;
        RECT 205.685 33.330 205.855 33.670 ;
        RECT 206.150 33.070 206.520 33.530 ;
        RECT 206.690 33.240 206.860 33.700 ;
        RECT 207.795 33.580 207.965 33.960 ;
        RECT 209.185 33.790 209.355 34.380 ;
        RECT 210.095 34.260 210.305 34.910 ;
        RECT 207.095 33.240 207.965 33.580 ;
        RECT 208.555 33.620 209.355 33.790 ;
        RECT 208.135 33.070 208.385 33.530 ;
        RECT 208.555 33.330 208.725 33.620 ;
        RECT 208.905 33.070 209.235 33.450 ;
        RECT 209.575 33.070 209.880 34.210 ;
        RECT 210.050 33.380 210.305 34.260 ;
        RECT 210.495 34.800 212.145 34.970 ;
        RECT 210.495 34.290 210.900 34.800 ;
        RECT 211.070 34.460 212.210 34.630 ;
        RECT 210.495 34.120 211.250 34.290 ;
        RECT 210.535 33.070 210.820 33.940 ;
        RECT 210.990 33.870 211.250 34.120 ;
        RECT 212.040 34.210 212.210 34.460 ;
        RECT 212.380 34.380 212.730 34.950 ;
        RECT 212.900 34.210 213.070 35.120 ;
        RECT 213.700 34.895 213.990 35.620 ;
        RECT 215.085 34.910 215.340 35.440 ;
        RECT 215.510 35.160 215.815 35.620 ;
        RECT 216.060 35.240 217.130 35.410 ;
        RECT 215.085 34.260 215.295 34.910 ;
        RECT 216.060 34.885 216.380 35.240 ;
        RECT 216.055 34.710 216.380 34.885 ;
        RECT 215.465 34.410 216.380 34.710 ;
        RECT 216.550 34.670 216.790 35.070 ;
        RECT 216.960 35.010 217.130 35.240 ;
        RECT 217.300 35.180 217.490 35.620 ;
        RECT 217.660 35.170 218.610 35.450 ;
        RECT 218.830 35.260 219.180 35.430 ;
        RECT 216.960 34.840 217.490 35.010 ;
        RECT 215.465 34.380 216.205 34.410 ;
        RECT 212.040 34.040 213.070 34.210 ;
        RECT 210.990 33.700 212.110 33.870 ;
        RECT 210.990 33.240 211.250 33.700 ;
        RECT 211.425 33.070 211.680 33.530 ;
        RECT 211.850 33.240 212.110 33.700 ;
        RECT 212.280 33.070 212.590 33.870 ;
        RECT 212.760 33.240 213.070 34.040 ;
        RECT 213.700 33.070 213.990 34.235 ;
        RECT 215.085 33.380 215.340 34.260 ;
        RECT 215.510 33.070 215.815 34.210 ;
        RECT 216.035 33.790 216.205 34.380 ;
        RECT 216.550 34.300 217.090 34.670 ;
        RECT 217.270 34.560 217.490 34.840 ;
        RECT 217.660 34.390 217.830 35.170 ;
        RECT 217.425 34.220 217.830 34.390 ;
        RECT 218.000 34.380 218.350 35.000 ;
        RECT 217.425 34.130 217.595 34.220 ;
        RECT 218.520 34.210 218.730 35.000 ;
        RECT 216.375 33.960 217.595 34.130 ;
        RECT 218.055 34.050 218.730 34.210 ;
        RECT 216.035 33.620 216.835 33.790 ;
        RECT 216.155 33.070 216.485 33.450 ;
        RECT 216.665 33.330 216.835 33.620 ;
        RECT 217.425 33.580 217.595 33.960 ;
        RECT 217.765 34.040 218.730 34.050 ;
        RECT 218.920 34.870 219.180 35.260 ;
        RECT 219.390 35.160 219.720 35.620 ;
        RECT 220.595 35.230 221.450 35.400 ;
        RECT 221.655 35.230 222.150 35.400 ;
        RECT 222.320 35.260 222.650 35.620 ;
        RECT 218.920 34.180 219.090 34.870 ;
        RECT 219.260 34.520 219.430 34.700 ;
        RECT 219.600 34.690 220.390 34.940 ;
        RECT 220.595 34.520 220.765 35.230 ;
        RECT 220.935 34.720 221.290 34.940 ;
        RECT 219.260 34.350 220.950 34.520 ;
        RECT 217.765 33.750 218.225 34.040 ;
        RECT 218.920 34.010 220.420 34.180 ;
        RECT 218.920 33.870 219.090 34.010 ;
        RECT 218.530 33.700 219.090 33.870 ;
        RECT 217.005 33.070 217.255 33.530 ;
        RECT 217.425 33.240 218.295 33.580 ;
        RECT 218.530 33.240 218.700 33.700 ;
        RECT 219.535 33.670 220.610 33.840 ;
        RECT 218.870 33.070 219.240 33.530 ;
        RECT 219.535 33.330 219.705 33.670 ;
        RECT 219.875 33.070 220.205 33.500 ;
        RECT 220.440 33.330 220.610 33.670 ;
        RECT 220.780 33.570 220.950 34.350 ;
        RECT 221.120 34.130 221.290 34.720 ;
        RECT 221.460 34.320 221.810 34.940 ;
        RECT 221.120 33.740 221.585 34.130 ;
        RECT 221.980 33.870 222.150 35.230 ;
        RECT 222.320 34.040 222.780 35.090 ;
        RECT 221.755 33.700 222.150 33.870 ;
        RECT 221.755 33.570 221.925 33.700 ;
        RECT 220.780 33.240 221.460 33.570 ;
        RECT 221.675 33.240 221.925 33.570 ;
        RECT 222.095 33.070 222.345 33.530 ;
        RECT 222.515 33.255 222.840 34.040 ;
        RECT 223.010 33.240 223.180 35.360 ;
        RECT 223.350 35.240 223.680 35.620 ;
        RECT 223.850 35.070 224.105 35.360 ;
        RECT 223.355 34.900 224.105 35.070 ;
        RECT 224.285 35.070 224.540 35.360 ;
        RECT 224.710 35.240 225.040 35.620 ;
        RECT 224.285 34.900 225.035 35.070 ;
        RECT 223.355 33.910 223.585 34.900 ;
        RECT 223.755 34.080 224.105 34.730 ;
        RECT 224.285 34.080 224.635 34.730 ;
        RECT 224.805 33.910 225.035 34.900 ;
        RECT 223.355 33.740 224.105 33.910 ;
        RECT 223.350 33.070 223.680 33.570 ;
        RECT 223.850 33.240 224.105 33.740 ;
        RECT 224.285 33.740 225.035 33.910 ;
        RECT 224.285 33.240 224.540 33.740 ;
        RECT 224.710 33.070 225.040 33.570 ;
        RECT 225.210 33.240 225.380 35.360 ;
        RECT 225.740 35.260 226.070 35.620 ;
        RECT 226.240 35.230 226.735 35.400 ;
        RECT 226.940 35.230 227.795 35.400 ;
        RECT 225.610 34.040 226.070 35.090 ;
        RECT 225.550 33.255 225.875 34.040 ;
        RECT 226.240 33.870 226.410 35.230 ;
        RECT 226.580 34.320 226.930 34.940 ;
        RECT 227.100 34.720 227.455 34.940 ;
        RECT 227.100 34.130 227.270 34.720 ;
        RECT 227.625 34.520 227.795 35.230 ;
        RECT 228.670 35.160 229.000 35.620 ;
        RECT 229.210 35.260 229.560 35.430 ;
        RECT 228.000 34.690 228.790 34.940 ;
        RECT 229.210 34.870 229.470 35.260 ;
        RECT 229.780 35.170 230.730 35.450 ;
        RECT 230.900 35.180 231.090 35.620 ;
        RECT 231.260 35.240 232.330 35.410 ;
        RECT 228.960 34.520 229.130 34.700 ;
        RECT 226.240 33.700 226.635 33.870 ;
        RECT 226.805 33.740 227.270 34.130 ;
        RECT 227.440 34.350 229.130 34.520 ;
        RECT 226.465 33.570 226.635 33.700 ;
        RECT 227.440 33.570 227.610 34.350 ;
        RECT 229.300 34.180 229.470 34.870 ;
        RECT 227.970 34.010 229.470 34.180 ;
        RECT 229.660 34.210 229.870 35.000 ;
        RECT 230.040 34.380 230.390 35.000 ;
        RECT 230.560 34.390 230.730 35.170 ;
        RECT 231.260 35.010 231.430 35.240 ;
        RECT 230.900 34.840 231.430 35.010 ;
        RECT 230.900 34.560 231.120 34.840 ;
        RECT 231.600 34.670 231.840 35.070 ;
        RECT 230.560 34.220 230.965 34.390 ;
        RECT 231.300 34.300 231.840 34.670 ;
        RECT 232.010 34.885 232.330 35.240 ;
        RECT 232.575 35.160 232.880 35.620 ;
        RECT 233.050 34.910 233.305 35.440 ;
        RECT 232.010 34.710 232.335 34.885 ;
        RECT 232.010 34.410 232.925 34.710 ;
        RECT 232.185 34.380 232.925 34.410 ;
        RECT 229.660 34.050 230.335 34.210 ;
        RECT 230.795 34.130 230.965 34.220 ;
        RECT 229.660 34.040 230.625 34.050 ;
        RECT 229.300 33.870 229.470 34.010 ;
        RECT 226.045 33.070 226.295 33.530 ;
        RECT 226.465 33.240 226.715 33.570 ;
        RECT 226.930 33.240 227.610 33.570 ;
        RECT 227.780 33.670 228.855 33.840 ;
        RECT 229.300 33.700 229.860 33.870 ;
        RECT 230.165 33.750 230.625 34.040 ;
        RECT 230.795 33.960 232.015 34.130 ;
        RECT 227.780 33.330 227.950 33.670 ;
        RECT 228.185 33.070 228.515 33.500 ;
        RECT 228.685 33.330 228.855 33.670 ;
        RECT 229.150 33.070 229.520 33.530 ;
        RECT 229.690 33.240 229.860 33.700 ;
        RECT 230.795 33.580 230.965 33.960 ;
        RECT 232.185 33.790 232.355 34.380 ;
        RECT 233.095 34.260 233.305 34.910 ;
        RECT 233.480 34.870 234.690 35.620 ;
        RECT 234.920 35.140 235.200 35.620 ;
        RECT 235.370 34.970 235.630 35.360 ;
        RECT 235.805 35.140 236.060 35.620 ;
        RECT 236.230 34.970 236.525 35.360 ;
        RECT 236.705 35.140 236.980 35.620 ;
        RECT 237.150 35.120 237.450 35.450 ;
        RECT 233.480 34.330 234.000 34.870 ;
        RECT 234.875 34.800 236.525 34.970 ;
        RECT 230.095 33.240 230.965 33.580 ;
        RECT 231.555 33.620 232.355 33.790 ;
        RECT 231.135 33.070 231.385 33.530 ;
        RECT 231.555 33.330 231.725 33.620 ;
        RECT 231.905 33.070 232.235 33.450 ;
        RECT 232.575 33.070 232.880 34.210 ;
        RECT 233.050 33.380 233.305 34.260 ;
        RECT 234.170 34.160 234.690 34.700 ;
        RECT 233.480 33.070 234.690 34.160 ;
        RECT 234.875 34.290 235.280 34.800 ;
        RECT 235.450 34.460 236.590 34.630 ;
        RECT 234.875 34.120 235.630 34.290 ;
        RECT 234.915 33.070 235.200 33.940 ;
        RECT 235.370 33.870 235.630 34.120 ;
        RECT 236.420 34.210 236.590 34.460 ;
        RECT 236.760 34.380 237.110 34.950 ;
        RECT 237.280 34.210 237.450 35.120 ;
        RECT 237.620 34.850 239.290 35.620 ;
        RECT 239.460 34.895 239.750 35.620 ;
        RECT 240.385 35.070 240.640 35.360 ;
        RECT 240.810 35.240 241.140 35.620 ;
        RECT 240.385 34.900 241.135 35.070 ;
        RECT 237.620 34.330 238.370 34.850 ;
        RECT 236.420 34.040 237.450 34.210 ;
        RECT 238.540 34.160 239.290 34.680 ;
        RECT 235.370 33.700 236.490 33.870 ;
        RECT 235.370 33.240 235.630 33.700 ;
        RECT 235.805 33.070 236.060 33.530 ;
        RECT 236.230 33.240 236.490 33.700 ;
        RECT 236.660 33.070 236.970 33.870 ;
        RECT 237.140 33.240 237.450 34.040 ;
        RECT 237.620 33.070 239.290 34.160 ;
        RECT 239.460 33.070 239.750 34.235 ;
        RECT 240.385 34.080 240.735 34.730 ;
        RECT 240.905 33.910 241.135 34.900 ;
        RECT 240.385 33.740 241.135 33.910 ;
        RECT 240.385 33.240 240.640 33.740 ;
        RECT 240.810 33.070 241.140 33.570 ;
        RECT 241.310 33.240 241.480 35.360 ;
        RECT 241.840 35.260 242.170 35.620 ;
        RECT 242.340 35.230 242.835 35.400 ;
        RECT 243.040 35.230 243.895 35.400 ;
        RECT 241.710 34.040 242.170 35.090 ;
        RECT 241.650 33.255 241.975 34.040 ;
        RECT 242.340 33.870 242.510 35.230 ;
        RECT 242.680 34.320 243.030 34.940 ;
        RECT 243.200 34.720 243.555 34.940 ;
        RECT 243.200 34.130 243.370 34.720 ;
        RECT 243.725 34.520 243.895 35.230 ;
        RECT 244.770 35.160 245.100 35.620 ;
        RECT 245.310 35.260 245.660 35.430 ;
        RECT 244.100 34.690 244.890 34.940 ;
        RECT 245.310 34.870 245.570 35.260 ;
        RECT 245.880 35.170 246.830 35.450 ;
        RECT 247.000 35.180 247.190 35.620 ;
        RECT 247.360 35.240 248.430 35.410 ;
        RECT 245.060 34.520 245.230 34.700 ;
        RECT 242.340 33.700 242.735 33.870 ;
        RECT 242.905 33.740 243.370 34.130 ;
        RECT 243.540 34.350 245.230 34.520 ;
        RECT 242.565 33.570 242.735 33.700 ;
        RECT 243.540 33.570 243.710 34.350 ;
        RECT 245.400 34.180 245.570 34.870 ;
        RECT 244.070 34.010 245.570 34.180 ;
        RECT 245.760 34.210 245.970 35.000 ;
        RECT 246.140 34.380 246.490 35.000 ;
        RECT 246.660 34.390 246.830 35.170 ;
        RECT 247.360 35.010 247.530 35.240 ;
        RECT 247.000 34.840 247.530 35.010 ;
        RECT 247.000 34.560 247.220 34.840 ;
        RECT 247.700 34.670 247.940 35.070 ;
        RECT 246.660 34.220 247.065 34.390 ;
        RECT 247.400 34.300 247.940 34.670 ;
        RECT 248.110 34.885 248.430 35.240 ;
        RECT 248.675 35.160 248.980 35.620 ;
        RECT 249.150 34.910 249.405 35.440 ;
        RECT 248.110 34.710 248.435 34.885 ;
        RECT 248.110 34.410 249.025 34.710 ;
        RECT 248.285 34.380 249.025 34.410 ;
        RECT 245.760 34.050 246.435 34.210 ;
        RECT 246.895 34.130 247.065 34.220 ;
        RECT 245.760 34.040 246.725 34.050 ;
        RECT 245.400 33.870 245.570 34.010 ;
        RECT 242.145 33.070 242.395 33.530 ;
        RECT 242.565 33.240 242.815 33.570 ;
        RECT 243.030 33.240 243.710 33.570 ;
        RECT 243.880 33.670 244.955 33.840 ;
        RECT 245.400 33.700 245.960 33.870 ;
        RECT 246.265 33.750 246.725 34.040 ;
        RECT 246.895 33.960 248.115 34.130 ;
        RECT 243.880 33.330 244.050 33.670 ;
        RECT 244.285 33.070 244.615 33.500 ;
        RECT 244.785 33.330 244.955 33.670 ;
        RECT 245.250 33.070 245.620 33.530 ;
        RECT 245.790 33.240 245.960 33.700 ;
        RECT 246.895 33.580 247.065 33.960 ;
        RECT 248.285 33.790 248.455 34.380 ;
        RECT 249.195 34.260 249.405 34.910 ;
        RECT 249.580 34.850 253.090 35.620 ;
        RECT 254.185 35.070 254.440 35.360 ;
        RECT 254.610 35.240 254.940 35.620 ;
        RECT 254.185 34.900 254.935 35.070 ;
        RECT 249.580 34.330 251.230 34.850 ;
        RECT 246.195 33.240 247.065 33.580 ;
        RECT 247.655 33.620 248.455 33.790 ;
        RECT 247.235 33.070 247.485 33.530 ;
        RECT 247.655 33.330 247.825 33.620 ;
        RECT 248.005 33.070 248.335 33.450 ;
        RECT 248.675 33.070 248.980 34.210 ;
        RECT 249.150 33.380 249.405 34.260 ;
        RECT 251.400 34.160 253.090 34.680 ;
        RECT 249.580 33.070 253.090 34.160 ;
        RECT 254.185 34.080 254.535 34.730 ;
        RECT 254.705 33.910 254.935 34.900 ;
        RECT 254.185 33.740 254.935 33.910 ;
        RECT 254.185 33.240 254.440 33.740 ;
        RECT 254.610 33.070 254.940 33.570 ;
        RECT 255.110 33.240 255.280 35.360 ;
        RECT 255.640 35.260 255.970 35.620 ;
        RECT 256.140 35.230 256.635 35.400 ;
        RECT 256.840 35.230 257.695 35.400 ;
        RECT 255.510 34.040 255.970 35.090 ;
        RECT 255.450 33.255 255.775 34.040 ;
        RECT 256.140 33.870 256.310 35.230 ;
        RECT 256.480 34.320 256.830 34.940 ;
        RECT 257.000 34.720 257.355 34.940 ;
        RECT 257.000 34.130 257.170 34.720 ;
        RECT 257.525 34.520 257.695 35.230 ;
        RECT 258.570 35.160 258.900 35.620 ;
        RECT 259.110 35.260 259.460 35.430 ;
        RECT 257.900 34.690 258.690 34.940 ;
        RECT 259.110 34.870 259.370 35.260 ;
        RECT 259.680 35.170 260.630 35.450 ;
        RECT 260.800 35.180 260.990 35.620 ;
        RECT 261.160 35.240 262.230 35.410 ;
        RECT 258.860 34.520 259.030 34.700 ;
        RECT 256.140 33.700 256.535 33.870 ;
        RECT 256.705 33.740 257.170 34.130 ;
        RECT 257.340 34.350 259.030 34.520 ;
        RECT 256.365 33.570 256.535 33.700 ;
        RECT 257.340 33.570 257.510 34.350 ;
        RECT 259.200 34.180 259.370 34.870 ;
        RECT 257.870 34.010 259.370 34.180 ;
        RECT 259.560 34.210 259.770 35.000 ;
        RECT 259.940 34.380 260.290 35.000 ;
        RECT 260.460 34.390 260.630 35.170 ;
        RECT 261.160 35.010 261.330 35.240 ;
        RECT 260.800 34.840 261.330 35.010 ;
        RECT 260.800 34.560 261.020 34.840 ;
        RECT 261.500 34.670 261.740 35.070 ;
        RECT 260.460 34.220 260.865 34.390 ;
        RECT 261.200 34.300 261.740 34.670 ;
        RECT 261.910 34.885 262.230 35.240 ;
        RECT 262.475 35.160 262.780 35.620 ;
        RECT 262.950 34.910 263.205 35.440 ;
        RECT 261.910 34.710 262.235 34.885 ;
        RECT 261.910 34.410 262.825 34.710 ;
        RECT 262.085 34.380 262.825 34.410 ;
        RECT 259.560 34.050 260.235 34.210 ;
        RECT 260.695 34.130 260.865 34.220 ;
        RECT 259.560 34.040 260.525 34.050 ;
        RECT 259.200 33.870 259.370 34.010 ;
        RECT 255.945 33.070 256.195 33.530 ;
        RECT 256.365 33.240 256.615 33.570 ;
        RECT 256.830 33.240 257.510 33.570 ;
        RECT 257.680 33.670 258.755 33.840 ;
        RECT 259.200 33.700 259.760 33.870 ;
        RECT 260.065 33.750 260.525 34.040 ;
        RECT 260.695 33.960 261.915 34.130 ;
        RECT 257.680 33.330 257.850 33.670 ;
        RECT 258.085 33.070 258.415 33.500 ;
        RECT 258.585 33.330 258.755 33.670 ;
        RECT 259.050 33.070 259.420 33.530 ;
        RECT 259.590 33.240 259.760 33.700 ;
        RECT 260.695 33.580 260.865 33.960 ;
        RECT 262.085 33.790 262.255 34.380 ;
        RECT 262.995 34.260 263.205 34.910 ;
        RECT 263.380 34.850 265.050 35.620 ;
        RECT 265.220 34.895 265.510 35.620 ;
        RECT 265.680 35.075 271.025 35.620 ;
        RECT 263.380 34.330 264.130 34.850 ;
        RECT 259.995 33.240 260.865 33.580 ;
        RECT 261.455 33.620 262.255 33.790 ;
        RECT 261.035 33.070 261.285 33.530 ;
        RECT 261.455 33.330 261.625 33.620 ;
        RECT 261.805 33.070 262.135 33.450 ;
        RECT 262.475 33.070 262.780 34.210 ;
        RECT 262.950 33.380 263.205 34.260 ;
        RECT 264.300 34.160 265.050 34.680 ;
        RECT 267.265 34.245 267.605 35.075 ;
        RECT 271.665 35.070 271.920 35.360 ;
        RECT 272.090 35.240 272.420 35.620 ;
        RECT 271.665 34.900 272.415 35.070 ;
        RECT 263.380 33.070 265.050 34.160 ;
        RECT 265.220 33.070 265.510 34.235 ;
        RECT 269.085 33.505 269.435 34.755 ;
        RECT 271.665 34.080 272.015 34.730 ;
        RECT 272.185 33.910 272.415 34.900 ;
        RECT 271.665 33.740 272.415 33.910 ;
        RECT 265.680 33.070 271.025 33.505 ;
        RECT 271.665 33.240 271.920 33.740 ;
        RECT 272.090 33.070 272.420 33.570 ;
        RECT 272.590 33.240 272.760 35.360 ;
        RECT 273.120 35.260 273.450 35.620 ;
        RECT 273.620 35.230 274.115 35.400 ;
        RECT 274.320 35.230 275.175 35.400 ;
        RECT 272.990 34.040 273.450 35.090 ;
        RECT 272.930 33.255 273.255 34.040 ;
        RECT 273.620 33.870 273.790 35.230 ;
        RECT 273.960 34.320 274.310 34.940 ;
        RECT 274.480 34.720 274.835 34.940 ;
        RECT 274.480 34.130 274.650 34.720 ;
        RECT 275.005 34.520 275.175 35.230 ;
        RECT 276.050 35.160 276.380 35.620 ;
        RECT 276.590 35.260 276.940 35.430 ;
        RECT 275.380 34.690 276.170 34.940 ;
        RECT 276.590 34.870 276.850 35.260 ;
        RECT 277.160 35.170 278.110 35.450 ;
        RECT 278.280 35.180 278.470 35.620 ;
        RECT 278.640 35.240 279.710 35.410 ;
        RECT 276.340 34.520 276.510 34.700 ;
        RECT 273.620 33.700 274.015 33.870 ;
        RECT 274.185 33.740 274.650 34.130 ;
        RECT 274.820 34.350 276.510 34.520 ;
        RECT 273.845 33.570 274.015 33.700 ;
        RECT 274.820 33.570 274.990 34.350 ;
        RECT 276.680 34.180 276.850 34.870 ;
        RECT 275.350 34.010 276.850 34.180 ;
        RECT 277.040 34.210 277.250 35.000 ;
        RECT 277.420 34.380 277.770 35.000 ;
        RECT 277.940 34.390 278.110 35.170 ;
        RECT 278.640 35.010 278.810 35.240 ;
        RECT 278.280 34.840 278.810 35.010 ;
        RECT 278.280 34.560 278.500 34.840 ;
        RECT 278.980 34.670 279.220 35.070 ;
        RECT 277.940 34.220 278.345 34.390 ;
        RECT 278.680 34.300 279.220 34.670 ;
        RECT 279.390 34.885 279.710 35.240 ;
        RECT 279.955 35.160 280.260 35.620 ;
        RECT 280.430 34.910 280.685 35.440 ;
        RECT 280.860 35.075 286.205 35.620 ;
        RECT 279.390 34.710 279.715 34.885 ;
        RECT 279.390 34.410 280.305 34.710 ;
        RECT 279.565 34.380 280.305 34.410 ;
        RECT 277.040 34.050 277.715 34.210 ;
        RECT 278.175 34.130 278.345 34.220 ;
        RECT 277.040 34.040 278.005 34.050 ;
        RECT 276.680 33.870 276.850 34.010 ;
        RECT 273.425 33.070 273.675 33.530 ;
        RECT 273.845 33.240 274.095 33.570 ;
        RECT 274.310 33.240 274.990 33.570 ;
        RECT 275.160 33.670 276.235 33.840 ;
        RECT 276.680 33.700 277.240 33.870 ;
        RECT 277.545 33.750 278.005 34.040 ;
        RECT 278.175 33.960 279.395 34.130 ;
        RECT 275.160 33.330 275.330 33.670 ;
        RECT 275.565 33.070 275.895 33.500 ;
        RECT 276.065 33.330 276.235 33.670 ;
        RECT 276.530 33.070 276.900 33.530 ;
        RECT 277.070 33.240 277.240 33.700 ;
        RECT 278.175 33.580 278.345 33.960 ;
        RECT 279.565 33.790 279.735 34.380 ;
        RECT 280.475 34.260 280.685 34.910 ;
        RECT 277.475 33.240 278.345 33.580 ;
        RECT 278.935 33.620 279.735 33.790 ;
        RECT 278.515 33.070 278.765 33.530 ;
        RECT 278.935 33.330 279.105 33.620 ;
        RECT 279.285 33.070 279.615 33.450 ;
        RECT 279.955 33.070 280.260 34.210 ;
        RECT 280.430 33.380 280.685 34.260 ;
        RECT 282.445 34.245 282.785 35.075 ;
        RECT 286.380 34.850 289.890 35.620 ;
        RECT 290.980 34.895 291.270 35.620 ;
        RECT 291.440 35.075 296.785 35.620 ;
        RECT 296.960 35.075 302.305 35.620 ;
        RECT 302.480 35.075 307.825 35.620 ;
        RECT 284.265 33.505 284.615 34.755 ;
        RECT 286.380 34.330 288.030 34.850 ;
        RECT 288.200 34.160 289.890 34.680 ;
        RECT 293.025 34.245 293.365 35.075 ;
        RECT 280.860 33.070 286.205 33.505 ;
        RECT 286.380 33.070 289.890 34.160 ;
        RECT 290.980 33.070 291.270 34.235 ;
        RECT 294.845 33.505 295.195 34.755 ;
        RECT 298.545 34.245 298.885 35.075 ;
        RECT 300.365 33.505 300.715 34.755 ;
        RECT 304.065 34.245 304.405 35.075 ;
        RECT 308.000 34.850 309.670 35.620 ;
        RECT 309.840 34.870 311.050 35.620 ;
        RECT 305.885 33.505 306.235 34.755 ;
        RECT 308.000 34.330 308.750 34.850 ;
        RECT 308.920 34.160 309.670 34.680 ;
        RECT 291.440 33.070 296.785 33.505 ;
        RECT 296.960 33.070 302.305 33.505 ;
        RECT 302.480 33.070 307.825 33.505 ;
        RECT 308.000 33.070 309.670 34.160 ;
        RECT 309.840 34.160 310.360 34.700 ;
        RECT 310.530 34.330 311.050 34.870 ;
        RECT 309.840 33.070 311.050 34.160 ;
        RECT 162.095 32.900 311.135 33.070 ;
        RECT 162.180 31.810 163.390 32.900 ;
        RECT 163.560 31.810 165.230 32.900 ;
        RECT 165.865 32.230 166.120 32.730 ;
        RECT 166.290 32.400 166.620 32.900 ;
        RECT 165.865 32.060 166.615 32.230 ;
        RECT 162.180 31.100 162.700 31.640 ;
        RECT 162.870 31.270 163.390 31.810 ;
        RECT 163.560 31.120 164.310 31.640 ;
        RECT 164.480 31.290 165.230 31.810 ;
        RECT 165.865 31.240 166.215 31.890 ;
        RECT 162.180 30.350 163.390 31.100 ;
        RECT 163.560 30.350 165.230 31.120 ;
        RECT 166.385 31.070 166.615 32.060 ;
        RECT 165.865 30.900 166.615 31.070 ;
        RECT 165.865 30.610 166.120 30.900 ;
        RECT 166.290 30.350 166.620 30.730 ;
        RECT 166.790 30.610 166.960 32.730 ;
        RECT 167.130 31.930 167.455 32.715 ;
        RECT 167.625 32.440 167.875 32.900 ;
        RECT 168.045 32.400 168.295 32.730 ;
        RECT 168.510 32.400 169.190 32.730 ;
        RECT 168.045 32.270 168.215 32.400 ;
        RECT 167.820 32.100 168.215 32.270 ;
        RECT 167.190 30.880 167.650 31.930 ;
        RECT 167.820 30.740 167.990 32.100 ;
        RECT 168.385 31.840 168.850 32.230 ;
        RECT 168.160 31.030 168.510 31.650 ;
        RECT 168.680 31.250 168.850 31.840 ;
        RECT 169.020 31.620 169.190 32.400 ;
        RECT 169.360 32.300 169.530 32.640 ;
        RECT 169.765 32.470 170.095 32.900 ;
        RECT 170.265 32.300 170.435 32.640 ;
        RECT 170.730 32.440 171.100 32.900 ;
        RECT 169.360 32.130 170.435 32.300 ;
        RECT 171.270 32.270 171.440 32.730 ;
        RECT 171.675 32.390 172.545 32.730 ;
        RECT 172.715 32.440 172.965 32.900 ;
        RECT 170.880 32.100 171.440 32.270 ;
        RECT 170.880 31.960 171.050 32.100 ;
        RECT 169.550 31.790 171.050 31.960 ;
        RECT 171.745 31.930 172.205 32.220 ;
        RECT 169.020 31.450 170.710 31.620 ;
        RECT 168.680 31.030 169.035 31.250 ;
        RECT 169.205 30.740 169.375 31.450 ;
        RECT 169.580 31.030 170.370 31.280 ;
        RECT 170.540 31.270 170.710 31.450 ;
        RECT 170.880 31.100 171.050 31.790 ;
        RECT 167.320 30.350 167.650 30.710 ;
        RECT 167.820 30.570 168.315 30.740 ;
        RECT 168.520 30.570 169.375 30.740 ;
        RECT 170.250 30.350 170.580 30.810 ;
        RECT 170.790 30.710 171.050 31.100 ;
        RECT 171.240 31.920 172.205 31.930 ;
        RECT 172.375 32.010 172.545 32.390 ;
        RECT 173.135 32.350 173.305 32.640 ;
        RECT 173.485 32.520 173.815 32.900 ;
        RECT 173.135 32.180 173.935 32.350 ;
        RECT 171.240 31.760 171.915 31.920 ;
        RECT 172.375 31.840 173.595 32.010 ;
        RECT 171.240 30.970 171.450 31.760 ;
        RECT 172.375 31.750 172.545 31.840 ;
        RECT 171.620 30.970 171.970 31.590 ;
        RECT 172.140 31.580 172.545 31.750 ;
        RECT 172.140 30.800 172.310 31.580 ;
        RECT 172.480 31.130 172.700 31.410 ;
        RECT 172.880 31.300 173.420 31.670 ;
        RECT 173.765 31.590 173.935 32.180 ;
        RECT 174.155 31.760 174.460 32.900 ;
        RECT 174.630 31.710 174.885 32.590 ;
        RECT 175.060 31.735 175.350 32.900 ;
        RECT 175.525 31.760 175.860 32.730 ;
        RECT 176.030 31.760 176.200 32.900 ;
        RECT 176.370 32.560 178.400 32.730 ;
        RECT 173.765 31.560 174.505 31.590 ;
        RECT 172.480 30.960 173.010 31.130 ;
        RECT 170.790 30.540 171.140 30.710 ;
        RECT 171.360 30.520 172.310 30.800 ;
        RECT 172.480 30.350 172.670 30.790 ;
        RECT 172.840 30.730 173.010 30.960 ;
        RECT 173.180 30.900 173.420 31.300 ;
        RECT 173.590 31.260 174.505 31.560 ;
        RECT 173.590 31.085 173.915 31.260 ;
        RECT 173.590 30.730 173.910 31.085 ;
        RECT 174.675 31.060 174.885 31.710 ;
        RECT 175.525 31.090 175.695 31.760 ;
        RECT 176.370 31.590 176.540 32.560 ;
        RECT 175.865 31.260 176.120 31.590 ;
        RECT 176.345 31.260 176.540 31.590 ;
        RECT 176.710 32.220 177.835 32.390 ;
        RECT 175.950 31.090 176.120 31.260 ;
        RECT 176.710 31.090 176.880 32.220 ;
        RECT 172.840 30.560 173.910 30.730 ;
        RECT 174.155 30.350 174.460 30.810 ;
        RECT 174.630 30.530 174.885 31.060 ;
        RECT 175.060 30.350 175.350 31.075 ;
        RECT 175.525 30.520 175.780 31.090 ;
        RECT 175.950 30.920 176.880 31.090 ;
        RECT 177.050 31.880 178.060 32.050 ;
        RECT 177.050 31.080 177.220 31.880 ;
        RECT 177.425 31.540 177.700 31.680 ;
        RECT 177.420 31.370 177.700 31.540 ;
        RECT 176.705 30.885 176.880 30.920 ;
        RECT 175.950 30.350 176.280 30.750 ;
        RECT 176.705 30.520 177.235 30.885 ;
        RECT 177.425 30.520 177.700 31.370 ;
        RECT 177.870 30.520 178.060 31.880 ;
        RECT 178.230 31.895 178.400 32.560 ;
        RECT 178.570 32.140 178.740 32.900 ;
        RECT 178.975 32.140 179.490 32.550 ;
        RECT 178.230 31.705 178.980 31.895 ;
        RECT 179.150 31.330 179.490 32.140 ;
        RECT 179.660 31.810 182.250 32.900 ;
        RECT 178.260 31.160 179.490 31.330 ;
        RECT 178.240 30.350 178.750 30.885 ;
        RECT 178.970 30.555 179.215 31.160 ;
        RECT 179.660 31.120 180.870 31.640 ;
        RECT 181.040 31.290 182.250 31.810 ;
        RECT 182.425 31.710 182.680 32.590 ;
        RECT 182.850 31.760 183.155 32.900 ;
        RECT 183.495 32.520 183.825 32.900 ;
        RECT 184.005 32.350 184.175 32.640 ;
        RECT 184.345 32.440 184.595 32.900 ;
        RECT 183.375 32.180 184.175 32.350 ;
        RECT 184.765 32.390 185.635 32.730 ;
        RECT 179.660 30.350 182.250 31.120 ;
        RECT 182.425 31.060 182.635 31.710 ;
        RECT 183.375 31.590 183.545 32.180 ;
        RECT 184.765 32.010 184.935 32.390 ;
        RECT 185.870 32.270 186.040 32.730 ;
        RECT 186.210 32.440 186.580 32.900 ;
        RECT 186.875 32.300 187.045 32.640 ;
        RECT 187.215 32.470 187.545 32.900 ;
        RECT 187.780 32.300 187.950 32.640 ;
        RECT 183.715 31.840 184.935 32.010 ;
        RECT 185.105 31.930 185.565 32.220 ;
        RECT 185.870 32.100 186.430 32.270 ;
        RECT 186.875 32.130 187.950 32.300 ;
        RECT 188.120 32.400 188.800 32.730 ;
        RECT 189.015 32.400 189.265 32.730 ;
        RECT 189.435 32.440 189.685 32.900 ;
        RECT 186.260 31.960 186.430 32.100 ;
        RECT 185.105 31.920 186.070 31.930 ;
        RECT 184.765 31.750 184.935 31.840 ;
        RECT 185.395 31.760 186.070 31.920 ;
        RECT 182.805 31.560 183.545 31.590 ;
        RECT 182.805 31.260 183.720 31.560 ;
        RECT 183.395 31.085 183.720 31.260 ;
        RECT 182.425 30.530 182.680 31.060 ;
        RECT 182.850 30.350 183.155 30.810 ;
        RECT 183.400 30.730 183.720 31.085 ;
        RECT 183.890 31.300 184.430 31.670 ;
        RECT 184.765 31.580 185.170 31.750 ;
        RECT 183.890 30.900 184.130 31.300 ;
        RECT 184.610 31.130 184.830 31.410 ;
        RECT 184.300 30.960 184.830 31.130 ;
        RECT 184.300 30.730 184.470 30.960 ;
        RECT 185.000 30.800 185.170 31.580 ;
        RECT 185.340 30.970 185.690 31.590 ;
        RECT 185.860 30.970 186.070 31.760 ;
        RECT 186.260 31.790 187.760 31.960 ;
        RECT 186.260 31.100 186.430 31.790 ;
        RECT 188.120 31.620 188.290 32.400 ;
        RECT 189.095 32.270 189.265 32.400 ;
        RECT 186.600 31.450 188.290 31.620 ;
        RECT 188.460 31.840 188.925 32.230 ;
        RECT 189.095 32.100 189.490 32.270 ;
        RECT 186.600 31.270 186.770 31.450 ;
        RECT 183.400 30.560 184.470 30.730 ;
        RECT 184.640 30.350 184.830 30.790 ;
        RECT 185.000 30.520 185.950 30.800 ;
        RECT 186.260 30.710 186.520 31.100 ;
        RECT 186.940 31.030 187.730 31.280 ;
        RECT 186.170 30.540 186.520 30.710 ;
        RECT 186.730 30.350 187.060 30.810 ;
        RECT 187.935 30.740 188.105 31.450 ;
        RECT 188.460 31.250 188.630 31.840 ;
        RECT 188.275 31.030 188.630 31.250 ;
        RECT 188.800 31.030 189.150 31.650 ;
        RECT 189.320 30.740 189.490 32.100 ;
        RECT 189.855 31.930 190.180 32.715 ;
        RECT 189.660 30.880 190.120 31.930 ;
        RECT 187.935 30.570 188.790 30.740 ;
        RECT 188.995 30.570 189.490 30.740 ;
        RECT 189.660 30.350 189.990 30.710 ;
        RECT 190.350 30.610 190.520 32.730 ;
        RECT 190.690 32.400 191.020 32.900 ;
        RECT 191.190 32.230 191.445 32.730 ;
        RECT 190.695 32.060 191.445 32.230 ;
        RECT 191.620 32.140 192.135 32.550 ;
        RECT 192.370 32.140 192.540 32.900 ;
        RECT 192.710 32.560 194.740 32.730 ;
        RECT 190.695 31.070 190.925 32.060 ;
        RECT 191.095 31.240 191.445 31.890 ;
        RECT 191.620 31.330 191.960 32.140 ;
        RECT 192.710 31.895 192.880 32.560 ;
        RECT 193.275 32.220 194.400 32.390 ;
        RECT 192.130 31.705 192.880 31.895 ;
        RECT 193.050 31.880 194.060 32.050 ;
        RECT 191.620 31.160 192.850 31.330 ;
        RECT 190.695 30.900 191.445 31.070 ;
        RECT 190.690 30.350 191.020 30.730 ;
        RECT 191.190 30.610 191.445 30.900 ;
        RECT 191.895 30.555 192.140 31.160 ;
        RECT 192.360 30.350 192.870 30.885 ;
        RECT 193.050 30.520 193.240 31.880 ;
        RECT 193.410 30.860 193.685 31.680 ;
        RECT 193.890 31.080 194.060 31.880 ;
        RECT 194.230 31.090 194.400 32.220 ;
        RECT 194.570 31.590 194.740 32.560 ;
        RECT 194.910 31.760 195.080 32.900 ;
        RECT 195.250 31.760 195.585 32.730 ;
        RECT 195.760 31.810 196.970 32.900 ;
        RECT 197.255 32.270 197.540 32.730 ;
        RECT 197.710 32.440 197.980 32.900 ;
        RECT 197.255 32.050 198.210 32.270 ;
        RECT 194.570 31.260 194.765 31.590 ;
        RECT 194.990 31.260 195.245 31.590 ;
        RECT 194.990 31.090 195.160 31.260 ;
        RECT 195.415 31.090 195.585 31.760 ;
        RECT 194.230 30.920 195.160 31.090 ;
        RECT 194.230 30.885 194.405 30.920 ;
        RECT 193.410 30.690 193.690 30.860 ;
        RECT 193.410 30.520 193.685 30.690 ;
        RECT 193.875 30.520 194.405 30.885 ;
        RECT 194.830 30.350 195.160 30.750 ;
        RECT 195.330 30.520 195.585 31.090 ;
        RECT 195.760 31.100 196.280 31.640 ;
        RECT 196.450 31.270 196.970 31.810 ;
        RECT 197.140 31.320 197.830 31.880 ;
        RECT 198.000 31.150 198.210 32.050 ;
        RECT 195.760 30.350 196.970 31.100 ;
        RECT 197.255 30.980 198.210 31.150 ;
        RECT 198.380 31.880 198.780 32.730 ;
        RECT 198.970 32.270 199.250 32.730 ;
        RECT 199.770 32.440 200.095 32.900 ;
        RECT 198.970 32.050 200.095 32.270 ;
        RECT 198.380 31.320 199.475 31.880 ;
        RECT 199.645 31.590 200.095 32.050 ;
        RECT 200.265 31.760 200.650 32.730 ;
        RECT 197.255 30.520 197.540 30.980 ;
        RECT 197.710 30.350 197.980 30.810 ;
        RECT 198.380 30.520 198.780 31.320 ;
        RECT 199.645 31.260 200.200 31.590 ;
        RECT 199.645 31.150 200.095 31.260 ;
        RECT 198.970 30.980 200.095 31.150 ;
        RECT 200.370 31.090 200.650 31.760 ;
        RECT 200.820 31.735 201.110 32.900 ;
        RECT 201.285 31.760 201.620 32.730 ;
        RECT 201.790 31.760 201.960 32.900 ;
        RECT 202.130 32.560 204.160 32.730 ;
        RECT 198.970 30.520 199.250 30.980 ;
        RECT 199.770 30.350 200.095 30.810 ;
        RECT 200.265 30.520 200.650 31.090 ;
        RECT 201.285 31.090 201.455 31.760 ;
        RECT 202.130 31.590 202.300 32.560 ;
        RECT 201.625 31.260 201.880 31.590 ;
        RECT 202.105 31.260 202.300 31.590 ;
        RECT 202.470 32.220 203.595 32.390 ;
        RECT 201.710 31.090 201.880 31.260 ;
        RECT 202.470 31.090 202.640 32.220 ;
        RECT 200.820 30.350 201.110 31.075 ;
        RECT 201.285 30.520 201.540 31.090 ;
        RECT 201.710 30.920 202.640 31.090 ;
        RECT 202.810 31.880 203.820 32.050 ;
        RECT 202.810 31.080 202.980 31.880 ;
        RECT 203.185 31.540 203.460 31.680 ;
        RECT 203.180 31.370 203.460 31.540 ;
        RECT 202.465 30.885 202.640 30.920 ;
        RECT 201.710 30.350 202.040 30.750 ;
        RECT 202.465 30.520 202.995 30.885 ;
        RECT 203.185 30.520 203.460 31.370 ;
        RECT 203.630 30.520 203.820 31.880 ;
        RECT 203.990 31.895 204.160 32.560 ;
        RECT 204.330 32.140 204.500 32.900 ;
        RECT 204.735 32.140 205.250 32.550 ;
        RECT 203.990 31.705 204.740 31.895 ;
        RECT 204.910 31.330 205.250 32.140 ;
        RECT 205.420 31.810 207.090 32.900 ;
        RECT 204.020 31.160 205.250 31.330 ;
        RECT 204.000 30.350 204.510 30.885 ;
        RECT 204.730 30.555 204.975 31.160 ;
        RECT 205.420 31.120 206.170 31.640 ;
        RECT 206.340 31.290 207.090 31.810 ;
        RECT 207.265 31.710 207.520 32.590 ;
        RECT 207.690 31.760 207.995 32.900 ;
        RECT 208.335 32.520 208.665 32.900 ;
        RECT 208.845 32.350 209.015 32.640 ;
        RECT 209.185 32.440 209.435 32.900 ;
        RECT 208.215 32.180 209.015 32.350 ;
        RECT 209.605 32.390 210.475 32.730 ;
        RECT 205.420 30.350 207.090 31.120 ;
        RECT 207.265 31.060 207.475 31.710 ;
        RECT 208.215 31.590 208.385 32.180 ;
        RECT 209.605 32.010 209.775 32.390 ;
        RECT 210.710 32.270 210.880 32.730 ;
        RECT 211.050 32.440 211.420 32.900 ;
        RECT 211.715 32.300 211.885 32.640 ;
        RECT 212.055 32.470 212.385 32.900 ;
        RECT 212.620 32.300 212.790 32.640 ;
        RECT 208.555 31.840 209.775 32.010 ;
        RECT 209.945 31.930 210.405 32.220 ;
        RECT 210.710 32.100 211.270 32.270 ;
        RECT 211.715 32.130 212.790 32.300 ;
        RECT 212.960 32.400 213.640 32.730 ;
        RECT 213.855 32.400 214.105 32.730 ;
        RECT 214.275 32.440 214.525 32.900 ;
        RECT 211.100 31.960 211.270 32.100 ;
        RECT 209.945 31.920 210.910 31.930 ;
        RECT 209.605 31.750 209.775 31.840 ;
        RECT 210.235 31.760 210.910 31.920 ;
        RECT 207.645 31.560 208.385 31.590 ;
        RECT 207.645 31.260 208.560 31.560 ;
        RECT 208.235 31.085 208.560 31.260 ;
        RECT 207.265 30.530 207.520 31.060 ;
        RECT 207.690 30.350 207.995 30.810 ;
        RECT 208.240 30.730 208.560 31.085 ;
        RECT 208.730 31.300 209.270 31.670 ;
        RECT 209.605 31.580 210.010 31.750 ;
        RECT 208.730 30.900 208.970 31.300 ;
        RECT 209.450 31.130 209.670 31.410 ;
        RECT 209.140 30.960 209.670 31.130 ;
        RECT 209.140 30.730 209.310 30.960 ;
        RECT 209.840 30.800 210.010 31.580 ;
        RECT 210.180 30.970 210.530 31.590 ;
        RECT 210.700 30.970 210.910 31.760 ;
        RECT 211.100 31.790 212.600 31.960 ;
        RECT 211.100 31.100 211.270 31.790 ;
        RECT 212.960 31.620 213.130 32.400 ;
        RECT 213.935 32.270 214.105 32.400 ;
        RECT 211.440 31.450 213.130 31.620 ;
        RECT 213.300 31.840 213.765 32.230 ;
        RECT 213.935 32.100 214.330 32.270 ;
        RECT 211.440 31.270 211.610 31.450 ;
        RECT 208.240 30.560 209.310 30.730 ;
        RECT 209.480 30.350 209.670 30.790 ;
        RECT 209.840 30.520 210.790 30.800 ;
        RECT 211.100 30.710 211.360 31.100 ;
        RECT 211.780 31.030 212.570 31.280 ;
        RECT 211.010 30.540 211.360 30.710 ;
        RECT 211.570 30.350 211.900 30.810 ;
        RECT 212.775 30.740 212.945 31.450 ;
        RECT 213.300 31.250 213.470 31.840 ;
        RECT 213.115 31.030 213.470 31.250 ;
        RECT 213.640 31.030 213.990 31.650 ;
        RECT 214.160 30.740 214.330 32.100 ;
        RECT 214.695 31.930 215.020 32.715 ;
        RECT 214.500 30.880 214.960 31.930 ;
        RECT 212.775 30.570 213.630 30.740 ;
        RECT 213.835 30.570 214.330 30.740 ;
        RECT 214.500 30.350 214.830 30.710 ;
        RECT 215.190 30.610 215.360 32.730 ;
        RECT 215.530 32.400 215.860 32.900 ;
        RECT 216.030 32.230 216.285 32.730 ;
        RECT 215.535 32.060 216.285 32.230 ;
        RECT 215.535 31.070 215.765 32.060 ;
        RECT 215.935 31.240 216.285 31.890 ;
        RECT 216.460 31.760 216.845 32.730 ;
        RECT 217.015 32.440 217.340 32.900 ;
        RECT 217.860 32.270 218.140 32.730 ;
        RECT 217.015 32.050 218.140 32.270 ;
        RECT 216.460 31.090 216.740 31.760 ;
        RECT 217.015 31.590 217.465 32.050 ;
        RECT 218.330 31.880 218.730 32.730 ;
        RECT 219.130 32.440 219.400 32.900 ;
        RECT 219.570 32.270 219.855 32.730 ;
        RECT 220.140 32.465 225.485 32.900 ;
        RECT 216.910 31.260 217.465 31.590 ;
        RECT 217.635 31.320 218.730 31.880 ;
        RECT 217.015 31.150 217.465 31.260 ;
        RECT 215.535 30.900 216.285 31.070 ;
        RECT 215.530 30.350 215.860 30.730 ;
        RECT 216.030 30.610 216.285 30.900 ;
        RECT 216.460 30.520 216.845 31.090 ;
        RECT 217.015 30.980 218.140 31.150 ;
        RECT 217.015 30.350 217.340 30.810 ;
        RECT 217.860 30.520 218.140 30.980 ;
        RECT 218.330 30.520 218.730 31.320 ;
        RECT 218.900 32.050 219.855 32.270 ;
        RECT 218.900 31.150 219.110 32.050 ;
        RECT 219.280 31.320 219.970 31.880 ;
        RECT 218.900 30.980 219.855 31.150 ;
        RECT 219.130 30.350 219.400 30.810 ;
        RECT 219.570 30.520 219.855 30.980 ;
        RECT 221.725 30.895 222.065 31.725 ;
        RECT 223.545 31.215 223.895 32.465 ;
        RECT 226.580 31.735 226.870 32.900 ;
        RECT 227.045 31.760 227.380 32.730 ;
        RECT 227.550 31.760 227.720 32.900 ;
        RECT 227.890 32.560 229.920 32.730 ;
        RECT 227.045 31.090 227.215 31.760 ;
        RECT 227.890 31.590 228.060 32.560 ;
        RECT 227.385 31.260 227.640 31.590 ;
        RECT 227.865 31.260 228.060 31.590 ;
        RECT 228.230 32.220 229.355 32.390 ;
        RECT 227.470 31.090 227.640 31.260 ;
        RECT 228.230 31.090 228.400 32.220 ;
        RECT 220.140 30.350 225.485 30.895 ;
        RECT 226.580 30.350 226.870 31.075 ;
        RECT 227.045 30.520 227.300 31.090 ;
        RECT 227.470 30.920 228.400 31.090 ;
        RECT 228.570 31.880 229.580 32.050 ;
        RECT 228.570 31.080 228.740 31.880 ;
        RECT 228.225 30.885 228.400 30.920 ;
        RECT 227.470 30.350 227.800 30.750 ;
        RECT 228.225 30.520 228.755 30.885 ;
        RECT 228.945 30.860 229.220 31.680 ;
        RECT 228.940 30.690 229.220 30.860 ;
        RECT 228.945 30.520 229.220 30.690 ;
        RECT 229.390 30.520 229.580 31.880 ;
        RECT 229.750 31.895 229.920 32.560 ;
        RECT 230.090 32.140 230.260 32.900 ;
        RECT 230.495 32.140 231.010 32.550 ;
        RECT 229.750 31.705 230.500 31.895 ;
        RECT 230.670 31.330 231.010 32.140 ;
        RECT 232.215 32.270 232.500 32.730 ;
        RECT 232.670 32.440 232.940 32.900 ;
        RECT 232.215 32.050 233.170 32.270 ;
        RECT 229.780 31.160 231.010 31.330 ;
        RECT 232.100 31.320 232.790 31.880 ;
        RECT 229.760 30.350 230.270 30.885 ;
        RECT 230.490 30.555 230.735 31.160 ;
        RECT 232.960 31.150 233.170 32.050 ;
        RECT 232.215 30.980 233.170 31.150 ;
        RECT 233.340 31.880 233.740 32.730 ;
        RECT 233.930 32.270 234.210 32.730 ;
        RECT 234.730 32.440 235.055 32.900 ;
        RECT 233.930 32.050 235.055 32.270 ;
        RECT 233.340 31.320 234.435 31.880 ;
        RECT 234.605 31.590 235.055 32.050 ;
        RECT 235.225 31.760 235.610 32.730 ;
        RECT 232.215 30.520 232.500 30.980 ;
        RECT 232.670 30.350 232.940 30.810 ;
        RECT 233.340 30.520 233.740 31.320 ;
        RECT 234.605 31.260 235.160 31.590 ;
        RECT 234.605 31.150 235.055 31.260 ;
        RECT 233.930 30.980 235.055 31.150 ;
        RECT 235.330 31.090 235.610 31.760 ;
        RECT 233.930 30.520 234.210 30.980 ;
        RECT 234.730 30.350 235.055 30.810 ;
        RECT 235.225 30.520 235.610 31.090 ;
        RECT 235.785 31.710 236.040 32.590 ;
        RECT 236.210 31.760 236.515 32.900 ;
        RECT 236.855 32.520 237.185 32.900 ;
        RECT 237.365 32.350 237.535 32.640 ;
        RECT 237.705 32.440 237.955 32.900 ;
        RECT 236.735 32.180 237.535 32.350 ;
        RECT 238.125 32.390 238.995 32.730 ;
        RECT 235.785 31.060 235.995 31.710 ;
        RECT 236.735 31.590 236.905 32.180 ;
        RECT 238.125 32.010 238.295 32.390 ;
        RECT 239.230 32.270 239.400 32.730 ;
        RECT 239.570 32.440 239.940 32.900 ;
        RECT 240.235 32.300 240.405 32.640 ;
        RECT 240.575 32.470 240.905 32.900 ;
        RECT 241.140 32.300 241.310 32.640 ;
        RECT 237.075 31.840 238.295 32.010 ;
        RECT 238.465 31.930 238.925 32.220 ;
        RECT 239.230 32.100 239.790 32.270 ;
        RECT 240.235 32.130 241.310 32.300 ;
        RECT 241.480 32.400 242.160 32.730 ;
        RECT 242.375 32.400 242.625 32.730 ;
        RECT 242.795 32.440 243.045 32.900 ;
        RECT 239.620 31.960 239.790 32.100 ;
        RECT 238.465 31.920 239.430 31.930 ;
        RECT 238.125 31.750 238.295 31.840 ;
        RECT 238.755 31.760 239.430 31.920 ;
        RECT 236.165 31.560 236.905 31.590 ;
        RECT 236.165 31.260 237.080 31.560 ;
        RECT 236.755 31.085 237.080 31.260 ;
        RECT 235.785 30.530 236.040 31.060 ;
        RECT 236.210 30.350 236.515 30.810 ;
        RECT 236.760 30.730 237.080 31.085 ;
        RECT 237.250 31.300 237.790 31.670 ;
        RECT 238.125 31.580 238.530 31.750 ;
        RECT 237.250 30.900 237.490 31.300 ;
        RECT 237.970 31.130 238.190 31.410 ;
        RECT 237.660 30.960 238.190 31.130 ;
        RECT 237.660 30.730 237.830 30.960 ;
        RECT 238.360 30.800 238.530 31.580 ;
        RECT 238.700 30.970 239.050 31.590 ;
        RECT 239.220 30.970 239.430 31.760 ;
        RECT 239.620 31.790 241.120 31.960 ;
        RECT 239.620 31.100 239.790 31.790 ;
        RECT 241.480 31.620 241.650 32.400 ;
        RECT 242.455 32.270 242.625 32.400 ;
        RECT 239.960 31.450 241.650 31.620 ;
        RECT 241.820 31.840 242.285 32.230 ;
        RECT 242.455 32.100 242.850 32.270 ;
        RECT 239.960 31.270 240.130 31.450 ;
        RECT 236.760 30.560 237.830 30.730 ;
        RECT 238.000 30.350 238.190 30.790 ;
        RECT 238.360 30.520 239.310 30.800 ;
        RECT 239.620 30.710 239.880 31.100 ;
        RECT 240.300 31.030 241.090 31.280 ;
        RECT 239.530 30.540 239.880 30.710 ;
        RECT 240.090 30.350 240.420 30.810 ;
        RECT 241.295 30.740 241.465 31.450 ;
        RECT 241.820 31.250 241.990 31.840 ;
        RECT 241.635 31.030 241.990 31.250 ;
        RECT 242.160 31.030 242.510 31.650 ;
        RECT 242.680 30.740 242.850 32.100 ;
        RECT 243.215 31.930 243.540 32.715 ;
        RECT 243.020 30.880 243.480 31.930 ;
        RECT 241.295 30.570 242.150 30.740 ;
        RECT 242.355 30.570 242.850 30.740 ;
        RECT 243.020 30.350 243.350 30.710 ;
        RECT 243.710 30.610 243.880 32.730 ;
        RECT 244.050 32.400 244.380 32.900 ;
        RECT 244.550 32.230 244.805 32.730 ;
        RECT 244.980 32.465 250.325 32.900 ;
        RECT 244.055 32.060 244.805 32.230 ;
        RECT 244.055 31.070 244.285 32.060 ;
        RECT 244.455 31.240 244.805 31.890 ;
        RECT 244.055 30.900 244.805 31.070 ;
        RECT 244.050 30.350 244.380 30.730 ;
        RECT 244.550 30.610 244.805 30.900 ;
        RECT 246.565 30.895 246.905 31.725 ;
        RECT 248.385 31.215 248.735 32.465 ;
        RECT 250.500 31.810 252.170 32.900 ;
        RECT 250.500 31.120 251.250 31.640 ;
        RECT 251.420 31.290 252.170 31.810 ;
        RECT 252.340 31.735 252.630 32.900 ;
        RECT 252.800 32.465 258.145 32.900 ;
        RECT 244.980 30.350 250.325 30.895 ;
        RECT 250.500 30.350 252.170 31.120 ;
        RECT 252.340 30.350 252.630 31.075 ;
        RECT 254.385 30.895 254.725 31.725 ;
        RECT 256.205 31.215 256.555 32.465 ;
        RECT 258.790 31.760 259.120 32.900 ;
        RECT 259.650 31.930 259.980 32.715 ;
        RECT 260.160 32.465 265.505 32.900 ;
        RECT 265.680 32.465 271.025 32.900 ;
        RECT 271.200 32.465 276.545 32.900 ;
        RECT 259.300 31.760 259.980 31.930 ;
        RECT 258.780 31.340 259.130 31.590 ;
        RECT 259.300 31.160 259.470 31.760 ;
        RECT 259.640 31.340 259.990 31.590 ;
        RECT 252.800 30.350 258.145 30.895 ;
        RECT 258.790 30.350 259.060 31.160 ;
        RECT 259.230 30.520 259.560 31.160 ;
        RECT 259.730 30.350 259.970 31.160 ;
        RECT 261.745 30.895 262.085 31.725 ;
        RECT 263.565 31.215 263.915 32.465 ;
        RECT 267.265 30.895 267.605 31.725 ;
        RECT 269.085 31.215 269.435 32.465 ;
        RECT 272.785 30.895 273.125 31.725 ;
        RECT 274.605 31.215 274.955 32.465 ;
        RECT 276.720 31.810 277.930 32.900 ;
        RECT 276.720 31.100 277.240 31.640 ;
        RECT 277.410 31.270 277.930 31.810 ;
        RECT 278.100 31.735 278.390 32.900 ;
        RECT 278.560 32.465 283.905 32.900 ;
        RECT 284.080 32.465 289.425 32.900 ;
        RECT 289.600 32.465 294.945 32.900 ;
        RECT 295.120 32.465 300.465 32.900 ;
        RECT 260.160 30.350 265.505 30.895 ;
        RECT 265.680 30.350 271.025 30.895 ;
        RECT 271.200 30.350 276.545 30.895 ;
        RECT 276.720 30.350 277.930 31.100 ;
        RECT 278.100 30.350 278.390 31.075 ;
        RECT 280.145 30.895 280.485 31.725 ;
        RECT 281.965 31.215 282.315 32.465 ;
        RECT 285.665 30.895 286.005 31.725 ;
        RECT 287.485 31.215 287.835 32.465 ;
        RECT 291.185 30.895 291.525 31.725 ;
        RECT 293.005 31.215 293.355 32.465 ;
        RECT 296.705 30.895 297.045 31.725 ;
        RECT 298.525 31.215 298.875 32.465 ;
        RECT 300.640 31.810 303.230 32.900 ;
        RECT 300.640 31.120 301.850 31.640 ;
        RECT 302.020 31.290 303.230 31.810 ;
        RECT 303.860 31.735 304.150 32.900 ;
        RECT 304.320 32.465 309.665 32.900 ;
        RECT 278.560 30.350 283.905 30.895 ;
        RECT 284.080 30.350 289.425 30.895 ;
        RECT 289.600 30.350 294.945 30.895 ;
        RECT 295.120 30.350 300.465 30.895 ;
        RECT 300.640 30.350 303.230 31.120 ;
        RECT 303.860 30.350 304.150 31.075 ;
        RECT 305.905 30.895 306.245 31.725 ;
        RECT 307.725 31.215 308.075 32.465 ;
        RECT 309.840 31.810 311.050 32.900 ;
        RECT 309.840 31.270 310.360 31.810 ;
        RECT 310.530 31.100 311.050 31.640 ;
        RECT 304.320 30.350 309.665 30.895 ;
        RECT 309.840 30.350 311.050 31.100 ;
        RECT 162.095 30.180 311.135 30.350 ;
        RECT 162.180 29.430 163.390 30.180 ;
        RECT 162.180 28.890 162.700 29.430 ;
        RECT 163.565 29.340 163.825 30.180 ;
        RECT 164.000 29.435 164.255 30.010 ;
        RECT 164.425 29.800 164.755 30.180 ;
        RECT 164.970 29.630 165.140 30.010 ;
        RECT 164.425 29.460 165.140 29.630 ;
        RECT 162.870 28.720 163.390 29.260 ;
        RECT 162.180 27.630 163.390 28.720 ;
        RECT 163.565 27.630 163.825 28.780 ;
        RECT 164.000 28.705 164.170 29.435 ;
        RECT 164.425 29.270 164.595 29.460 ;
        RECT 165.400 29.410 167.990 30.180 ;
        RECT 168.620 29.440 169.005 30.010 ;
        RECT 169.175 29.720 169.500 30.180 ;
        RECT 170.020 29.550 170.300 30.010 ;
        RECT 164.340 28.940 164.595 29.270 ;
        RECT 164.425 28.730 164.595 28.940 ;
        RECT 164.875 28.910 165.230 29.280 ;
        RECT 165.400 28.890 166.610 29.410 ;
        RECT 164.000 27.800 164.255 28.705 ;
        RECT 164.425 28.560 165.140 28.730 ;
        RECT 166.780 28.720 167.990 29.240 ;
        RECT 164.425 27.630 164.755 28.390 ;
        RECT 164.970 27.800 165.140 28.560 ;
        RECT 165.400 27.630 167.990 28.720 ;
        RECT 168.620 28.770 168.900 29.440 ;
        RECT 169.175 29.380 170.300 29.550 ;
        RECT 169.175 29.270 169.625 29.380 ;
        RECT 169.070 28.940 169.625 29.270 ;
        RECT 170.490 29.210 170.890 30.010 ;
        RECT 171.290 29.720 171.560 30.180 ;
        RECT 171.730 29.550 172.015 30.010 ;
        RECT 168.620 27.800 169.005 28.770 ;
        RECT 169.175 28.480 169.625 28.940 ;
        RECT 169.795 28.650 170.890 29.210 ;
        RECT 169.175 28.260 170.300 28.480 ;
        RECT 169.175 27.630 169.500 28.090 ;
        RECT 170.020 27.800 170.300 28.260 ;
        RECT 170.490 27.800 170.890 28.650 ;
        RECT 171.060 29.380 172.015 29.550 ;
        RECT 172.305 29.440 172.560 30.010 ;
        RECT 172.730 29.780 173.060 30.180 ;
        RECT 173.485 29.645 174.015 30.010 ;
        RECT 173.485 29.610 173.660 29.645 ;
        RECT 172.730 29.440 173.660 29.610 ;
        RECT 174.205 29.500 174.480 30.010 ;
        RECT 171.060 28.480 171.270 29.380 ;
        RECT 171.440 28.650 172.130 29.210 ;
        RECT 172.305 28.770 172.475 29.440 ;
        RECT 172.730 29.270 172.900 29.440 ;
        RECT 172.645 28.940 172.900 29.270 ;
        RECT 173.125 28.940 173.320 29.270 ;
        RECT 171.060 28.260 172.015 28.480 ;
        RECT 171.290 27.630 171.560 28.090 ;
        RECT 171.730 27.800 172.015 28.260 ;
        RECT 172.305 27.800 172.640 28.770 ;
        RECT 172.810 27.630 172.980 28.770 ;
        RECT 173.150 27.970 173.320 28.940 ;
        RECT 173.490 28.310 173.660 29.440 ;
        RECT 173.830 28.650 174.000 29.450 ;
        RECT 174.200 29.330 174.480 29.500 ;
        RECT 174.205 28.850 174.480 29.330 ;
        RECT 174.650 28.650 174.840 30.010 ;
        RECT 175.020 29.645 175.530 30.180 ;
        RECT 175.750 29.370 175.995 29.975 ;
        RECT 176.555 29.550 176.840 30.010 ;
        RECT 177.010 29.720 177.280 30.180 ;
        RECT 176.555 29.380 177.510 29.550 ;
        RECT 175.040 29.200 176.270 29.370 ;
        RECT 173.830 28.480 174.840 28.650 ;
        RECT 175.010 28.635 175.760 28.825 ;
        RECT 173.490 28.140 174.615 28.310 ;
        RECT 175.010 27.970 175.180 28.635 ;
        RECT 175.930 28.390 176.270 29.200 ;
        RECT 176.440 28.650 177.130 29.210 ;
        RECT 177.300 28.480 177.510 29.380 ;
        RECT 173.150 27.800 175.180 27.970 ;
        RECT 175.350 27.630 175.520 28.390 ;
        RECT 175.755 27.980 176.270 28.390 ;
        RECT 176.555 28.260 177.510 28.480 ;
        RECT 177.680 29.210 178.080 30.010 ;
        RECT 178.270 29.550 178.550 30.010 ;
        RECT 179.070 29.720 179.395 30.180 ;
        RECT 178.270 29.380 179.395 29.550 ;
        RECT 179.565 29.440 179.950 30.010 ;
        RECT 178.945 29.270 179.395 29.380 ;
        RECT 177.680 28.650 178.775 29.210 ;
        RECT 178.945 28.940 179.500 29.270 ;
        RECT 176.555 27.800 176.840 28.260 ;
        RECT 177.010 27.630 177.280 28.090 ;
        RECT 177.680 27.800 178.080 28.650 ;
        RECT 178.945 28.480 179.395 28.940 ;
        RECT 179.670 28.770 179.950 29.440 ;
        RECT 180.235 29.550 180.520 30.010 ;
        RECT 180.690 29.720 180.960 30.180 ;
        RECT 180.235 29.380 181.190 29.550 ;
        RECT 178.270 28.260 179.395 28.480 ;
        RECT 178.270 27.800 178.550 28.260 ;
        RECT 179.070 27.630 179.395 28.090 ;
        RECT 179.565 27.800 179.950 28.770 ;
        RECT 180.120 28.650 180.810 29.210 ;
        RECT 180.980 28.480 181.190 29.380 ;
        RECT 180.235 28.260 181.190 28.480 ;
        RECT 181.360 29.210 181.760 30.010 ;
        RECT 181.950 29.550 182.230 30.010 ;
        RECT 182.750 29.720 183.075 30.180 ;
        RECT 181.950 29.380 183.075 29.550 ;
        RECT 183.245 29.440 183.630 30.010 ;
        RECT 182.625 29.270 183.075 29.380 ;
        RECT 181.360 28.650 182.455 29.210 ;
        RECT 182.625 28.940 183.180 29.270 ;
        RECT 180.235 27.800 180.520 28.260 ;
        RECT 180.690 27.630 180.960 28.090 ;
        RECT 181.360 27.800 181.760 28.650 ;
        RECT 182.625 28.480 183.075 28.940 ;
        RECT 183.350 28.770 183.630 29.440 ;
        RECT 181.950 28.260 183.075 28.480 ;
        RECT 181.950 27.800 182.230 28.260 ;
        RECT 182.750 27.630 183.075 28.090 ;
        RECT 183.245 27.800 183.630 28.770 ;
        RECT 183.805 29.440 184.060 30.010 ;
        RECT 184.230 29.780 184.560 30.180 ;
        RECT 184.985 29.645 185.515 30.010 ;
        RECT 184.985 29.610 185.160 29.645 ;
        RECT 184.230 29.440 185.160 29.610 ;
        RECT 185.705 29.500 185.980 30.010 ;
        RECT 183.805 28.770 183.975 29.440 ;
        RECT 184.230 29.270 184.400 29.440 ;
        RECT 184.145 28.940 184.400 29.270 ;
        RECT 184.625 28.940 184.820 29.270 ;
        RECT 183.805 27.800 184.140 28.770 ;
        RECT 184.310 27.630 184.480 28.770 ;
        RECT 184.650 27.970 184.820 28.940 ;
        RECT 184.990 28.310 185.160 29.440 ;
        RECT 185.330 28.650 185.500 29.450 ;
        RECT 185.700 29.330 185.980 29.500 ;
        RECT 185.705 28.850 185.980 29.330 ;
        RECT 186.150 28.650 186.340 30.010 ;
        RECT 186.520 29.645 187.030 30.180 ;
        RECT 187.250 29.370 187.495 29.975 ;
        RECT 187.940 29.455 188.230 30.180 ;
        RECT 188.405 29.440 188.660 30.010 ;
        RECT 188.830 29.780 189.160 30.180 ;
        RECT 189.585 29.645 190.115 30.010 ;
        RECT 189.585 29.610 189.760 29.645 ;
        RECT 188.830 29.440 189.760 29.610 ;
        RECT 186.540 29.200 187.770 29.370 ;
        RECT 185.330 28.480 186.340 28.650 ;
        RECT 186.510 28.635 187.260 28.825 ;
        RECT 184.990 28.140 186.115 28.310 ;
        RECT 186.510 27.970 186.680 28.635 ;
        RECT 187.430 28.390 187.770 29.200 ;
        RECT 184.650 27.800 186.680 27.970 ;
        RECT 186.850 27.630 187.020 28.390 ;
        RECT 187.255 27.980 187.770 28.390 ;
        RECT 187.940 27.630 188.230 28.795 ;
        RECT 188.405 28.770 188.575 29.440 ;
        RECT 188.830 29.270 189.000 29.440 ;
        RECT 188.745 28.940 189.000 29.270 ;
        RECT 189.225 28.940 189.420 29.270 ;
        RECT 188.405 27.800 188.740 28.770 ;
        RECT 188.910 27.630 189.080 28.770 ;
        RECT 189.250 27.970 189.420 28.940 ;
        RECT 189.590 28.310 189.760 29.440 ;
        RECT 189.930 28.650 190.100 29.450 ;
        RECT 190.305 29.160 190.580 30.010 ;
        RECT 190.300 28.990 190.580 29.160 ;
        RECT 190.305 28.850 190.580 28.990 ;
        RECT 190.750 28.650 190.940 30.010 ;
        RECT 191.120 29.645 191.630 30.180 ;
        RECT 191.850 29.370 192.095 29.975 ;
        RECT 193.000 29.440 193.385 30.010 ;
        RECT 193.555 29.720 193.880 30.180 ;
        RECT 194.400 29.550 194.680 30.010 ;
        RECT 191.140 29.200 192.370 29.370 ;
        RECT 189.930 28.480 190.940 28.650 ;
        RECT 191.110 28.635 191.860 28.825 ;
        RECT 189.590 28.140 190.715 28.310 ;
        RECT 191.110 27.970 191.280 28.635 ;
        RECT 192.030 28.390 192.370 29.200 ;
        RECT 189.250 27.800 191.280 27.970 ;
        RECT 191.450 27.630 191.620 28.390 ;
        RECT 191.855 27.980 192.370 28.390 ;
        RECT 193.000 28.770 193.280 29.440 ;
        RECT 193.555 29.380 194.680 29.550 ;
        RECT 193.555 29.270 194.005 29.380 ;
        RECT 193.450 28.940 194.005 29.270 ;
        RECT 194.870 29.210 195.270 30.010 ;
        RECT 195.670 29.720 195.940 30.180 ;
        RECT 196.110 29.550 196.395 30.010 ;
        RECT 193.000 27.800 193.385 28.770 ;
        RECT 193.555 28.480 194.005 28.940 ;
        RECT 194.175 28.650 195.270 29.210 ;
        RECT 193.555 28.260 194.680 28.480 ;
        RECT 193.555 27.630 193.880 28.090 ;
        RECT 194.400 27.800 194.680 28.260 ;
        RECT 194.870 27.800 195.270 28.650 ;
        RECT 195.440 29.380 196.395 29.550 ;
        RECT 196.685 29.470 196.940 30.000 ;
        RECT 197.110 29.720 197.415 30.180 ;
        RECT 197.660 29.800 198.730 29.970 ;
        RECT 195.440 28.480 195.650 29.380 ;
        RECT 195.820 28.650 196.510 29.210 ;
        RECT 196.685 28.820 196.895 29.470 ;
        RECT 197.660 29.445 197.980 29.800 ;
        RECT 197.655 29.270 197.980 29.445 ;
        RECT 197.065 28.970 197.980 29.270 ;
        RECT 198.150 29.230 198.390 29.630 ;
        RECT 198.560 29.570 198.730 29.800 ;
        RECT 198.900 29.740 199.090 30.180 ;
        RECT 199.260 29.730 200.210 30.010 ;
        RECT 200.430 29.820 200.780 29.990 ;
        RECT 198.560 29.400 199.090 29.570 ;
        RECT 197.065 28.940 197.805 28.970 ;
        RECT 195.440 28.260 196.395 28.480 ;
        RECT 195.670 27.630 195.940 28.090 ;
        RECT 196.110 27.800 196.395 28.260 ;
        RECT 196.685 27.940 196.940 28.820 ;
        RECT 197.110 27.630 197.415 28.770 ;
        RECT 197.635 28.350 197.805 28.940 ;
        RECT 198.150 28.860 198.690 29.230 ;
        RECT 198.870 29.120 199.090 29.400 ;
        RECT 199.260 28.950 199.430 29.730 ;
        RECT 199.025 28.780 199.430 28.950 ;
        RECT 199.600 28.940 199.950 29.560 ;
        RECT 199.025 28.690 199.195 28.780 ;
        RECT 200.120 28.770 200.330 29.560 ;
        RECT 197.975 28.520 199.195 28.690 ;
        RECT 199.655 28.610 200.330 28.770 ;
        RECT 197.635 28.180 198.435 28.350 ;
        RECT 197.755 27.630 198.085 28.010 ;
        RECT 198.265 27.890 198.435 28.180 ;
        RECT 199.025 28.140 199.195 28.520 ;
        RECT 199.365 28.600 200.330 28.610 ;
        RECT 200.520 29.430 200.780 29.820 ;
        RECT 200.990 29.720 201.320 30.180 ;
        RECT 202.195 29.790 203.050 29.960 ;
        RECT 203.255 29.790 203.750 29.960 ;
        RECT 203.920 29.820 204.250 30.180 ;
        RECT 200.520 28.740 200.690 29.430 ;
        RECT 200.860 29.080 201.030 29.260 ;
        RECT 201.200 29.250 201.990 29.500 ;
        RECT 202.195 29.080 202.365 29.790 ;
        RECT 202.535 29.280 202.890 29.500 ;
        RECT 200.860 28.910 202.550 29.080 ;
        RECT 199.365 28.310 199.825 28.600 ;
        RECT 200.520 28.570 202.020 28.740 ;
        RECT 200.520 28.430 200.690 28.570 ;
        RECT 200.130 28.260 200.690 28.430 ;
        RECT 198.605 27.630 198.855 28.090 ;
        RECT 199.025 27.800 199.895 28.140 ;
        RECT 200.130 27.800 200.300 28.260 ;
        RECT 201.135 28.230 202.210 28.400 ;
        RECT 200.470 27.630 200.840 28.090 ;
        RECT 201.135 27.890 201.305 28.230 ;
        RECT 201.475 27.630 201.805 28.060 ;
        RECT 202.040 27.890 202.210 28.230 ;
        RECT 202.380 28.130 202.550 28.910 ;
        RECT 202.720 28.690 202.890 29.280 ;
        RECT 203.060 28.880 203.410 29.500 ;
        RECT 202.720 28.300 203.185 28.690 ;
        RECT 203.580 28.430 203.750 29.790 ;
        RECT 203.920 28.600 204.380 29.650 ;
        RECT 203.355 28.260 203.750 28.430 ;
        RECT 203.355 28.130 203.525 28.260 ;
        RECT 202.380 27.800 203.060 28.130 ;
        RECT 203.275 27.800 203.525 28.130 ;
        RECT 203.695 27.630 203.945 28.090 ;
        RECT 204.115 27.815 204.440 28.600 ;
        RECT 204.610 27.800 204.780 29.920 ;
        RECT 204.950 29.800 205.280 30.180 ;
        RECT 205.450 29.630 205.705 29.920 ;
        RECT 204.955 29.460 205.705 29.630 ;
        RECT 204.955 28.470 205.185 29.460 ;
        RECT 205.880 29.410 208.470 30.180 ;
        RECT 208.640 29.440 209.025 30.010 ;
        RECT 209.195 29.720 209.520 30.180 ;
        RECT 210.040 29.550 210.320 30.010 ;
        RECT 205.355 28.640 205.705 29.290 ;
        RECT 205.880 28.890 207.090 29.410 ;
        RECT 207.260 28.720 208.470 29.240 ;
        RECT 204.955 28.300 205.705 28.470 ;
        RECT 204.950 27.630 205.280 28.130 ;
        RECT 205.450 27.800 205.705 28.300 ;
        RECT 205.880 27.630 208.470 28.720 ;
        RECT 208.640 28.770 208.920 29.440 ;
        RECT 209.195 29.380 210.320 29.550 ;
        RECT 209.195 29.270 209.645 29.380 ;
        RECT 209.090 28.940 209.645 29.270 ;
        RECT 210.510 29.210 210.910 30.010 ;
        RECT 211.310 29.720 211.580 30.180 ;
        RECT 211.750 29.550 212.035 30.010 ;
        RECT 208.640 27.800 209.025 28.770 ;
        RECT 209.195 28.480 209.645 28.940 ;
        RECT 209.815 28.650 210.910 29.210 ;
        RECT 209.195 28.260 210.320 28.480 ;
        RECT 209.195 27.630 209.520 28.090 ;
        RECT 210.040 27.800 210.320 28.260 ;
        RECT 210.510 27.800 210.910 28.650 ;
        RECT 211.080 29.380 212.035 29.550 ;
        RECT 212.320 29.430 213.530 30.180 ;
        RECT 213.700 29.455 213.990 30.180 ;
        RECT 214.160 29.635 219.505 30.180 ;
        RECT 219.680 29.635 225.025 30.180 ;
        RECT 225.200 29.635 230.545 30.180 ;
        RECT 230.720 29.635 236.065 30.180 ;
        RECT 211.080 28.480 211.290 29.380 ;
        RECT 211.460 28.650 212.150 29.210 ;
        RECT 212.320 28.890 212.840 29.430 ;
        RECT 213.010 28.720 213.530 29.260 ;
        RECT 215.745 28.805 216.085 29.635 ;
        RECT 211.080 28.260 212.035 28.480 ;
        RECT 211.310 27.630 211.580 28.090 ;
        RECT 211.750 27.800 212.035 28.260 ;
        RECT 212.320 27.630 213.530 28.720 ;
        RECT 213.700 27.630 213.990 28.795 ;
        RECT 217.565 28.065 217.915 29.315 ;
        RECT 221.265 28.805 221.605 29.635 ;
        RECT 223.085 28.065 223.435 29.315 ;
        RECT 226.785 28.805 227.125 29.635 ;
        RECT 228.605 28.065 228.955 29.315 ;
        RECT 232.305 28.805 232.645 29.635 ;
        RECT 236.240 29.410 238.830 30.180 ;
        RECT 239.460 29.455 239.750 30.180 ;
        RECT 239.920 29.635 245.265 30.180 ;
        RECT 245.440 29.635 250.785 30.180 ;
        RECT 250.960 29.635 256.305 30.180 ;
        RECT 256.480 29.635 261.825 30.180 ;
        RECT 234.125 28.065 234.475 29.315 ;
        RECT 236.240 28.890 237.450 29.410 ;
        RECT 237.620 28.720 238.830 29.240 ;
        RECT 241.505 28.805 241.845 29.635 ;
        RECT 214.160 27.630 219.505 28.065 ;
        RECT 219.680 27.630 225.025 28.065 ;
        RECT 225.200 27.630 230.545 28.065 ;
        RECT 230.720 27.630 236.065 28.065 ;
        RECT 236.240 27.630 238.830 28.720 ;
        RECT 239.460 27.630 239.750 28.795 ;
        RECT 243.325 28.065 243.675 29.315 ;
        RECT 247.025 28.805 247.365 29.635 ;
        RECT 248.845 28.065 249.195 29.315 ;
        RECT 252.545 28.805 252.885 29.635 ;
        RECT 254.365 28.065 254.715 29.315 ;
        RECT 258.065 28.805 258.405 29.635 ;
        RECT 262.000 29.410 264.590 30.180 ;
        RECT 265.220 29.455 265.510 30.180 ;
        RECT 265.680 29.635 271.025 30.180 ;
        RECT 271.200 29.635 276.545 30.180 ;
        RECT 276.720 29.635 282.065 30.180 ;
        RECT 282.240 29.635 287.585 30.180 ;
        RECT 259.885 28.065 260.235 29.315 ;
        RECT 262.000 28.890 263.210 29.410 ;
        RECT 263.380 28.720 264.590 29.240 ;
        RECT 267.265 28.805 267.605 29.635 ;
        RECT 239.920 27.630 245.265 28.065 ;
        RECT 245.440 27.630 250.785 28.065 ;
        RECT 250.960 27.630 256.305 28.065 ;
        RECT 256.480 27.630 261.825 28.065 ;
        RECT 262.000 27.630 264.590 28.720 ;
        RECT 265.220 27.630 265.510 28.795 ;
        RECT 269.085 28.065 269.435 29.315 ;
        RECT 272.785 28.805 273.125 29.635 ;
        RECT 274.605 28.065 274.955 29.315 ;
        RECT 278.305 28.805 278.645 29.635 ;
        RECT 280.125 28.065 280.475 29.315 ;
        RECT 283.825 28.805 284.165 29.635 ;
        RECT 287.760 29.410 290.350 30.180 ;
        RECT 290.980 29.455 291.270 30.180 ;
        RECT 291.440 29.635 296.785 30.180 ;
        RECT 296.960 29.635 302.305 30.180 ;
        RECT 302.480 29.635 307.825 30.180 ;
        RECT 285.645 28.065 285.995 29.315 ;
        RECT 287.760 28.890 288.970 29.410 ;
        RECT 289.140 28.720 290.350 29.240 ;
        RECT 293.025 28.805 293.365 29.635 ;
        RECT 265.680 27.630 271.025 28.065 ;
        RECT 271.200 27.630 276.545 28.065 ;
        RECT 276.720 27.630 282.065 28.065 ;
        RECT 282.240 27.630 287.585 28.065 ;
        RECT 287.760 27.630 290.350 28.720 ;
        RECT 290.980 27.630 291.270 28.795 ;
        RECT 294.845 28.065 295.195 29.315 ;
        RECT 298.545 28.805 298.885 29.635 ;
        RECT 300.365 28.065 300.715 29.315 ;
        RECT 304.065 28.805 304.405 29.635 ;
        RECT 308.000 29.410 309.670 30.180 ;
        RECT 309.840 29.430 311.050 30.180 ;
        RECT 305.885 28.065 306.235 29.315 ;
        RECT 308.000 28.890 308.750 29.410 ;
        RECT 308.920 28.720 309.670 29.240 ;
        RECT 291.440 27.630 296.785 28.065 ;
        RECT 296.960 27.630 302.305 28.065 ;
        RECT 302.480 27.630 307.825 28.065 ;
        RECT 308.000 27.630 309.670 28.720 ;
        RECT 309.840 28.720 310.360 29.260 ;
        RECT 310.530 28.890 311.050 29.430 ;
        RECT 309.840 27.630 311.050 28.720 ;
        RECT 162.095 27.460 311.135 27.630 ;
        RECT 162.180 26.370 163.390 27.460 ;
        RECT 163.560 27.025 168.905 27.460 ;
        RECT 162.180 25.660 162.700 26.200 ;
        RECT 162.870 25.830 163.390 26.370 ;
        RECT 162.180 24.910 163.390 25.660 ;
        RECT 165.145 25.455 165.485 26.285 ;
        RECT 166.965 25.775 167.315 27.025 ;
        RECT 169.080 26.370 170.750 27.460 ;
        RECT 169.080 25.680 169.830 26.200 ;
        RECT 170.000 25.850 170.750 26.370 ;
        RECT 171.380 26.320 171.765 27.290 ;
        RECT 171.935 27.000 172.260 27.460 ;
        RECT 172.780 26.830 173.060 27.290 ;
        RECT 171.935 26.610 173.060 26.830 ;
        RECT 163.560 24.910 168.905 25.455 ;
        RECT 169.080 24.910 170.750 25.680 ;
        RECT 171.380 25.650 171.660 26.320 ;
        RECT 171.935 26.150 172.385 26.610 ;
        RECT 173.250 26.440 173.650 27.290 ;
        RECT 174.050 27.000 174.320 27.460 ;
        RECT 174.490 26.830 174.775 27.290 ;
        RECT 171.830 25.820 172.385 26.150 ;
        RECT 172.555 25.880 173.650 26.440 ;
        RECT 171.935 25.710 172.385 25.820 ;
        RECT 171.380 25.080 171.765 25.650 ;
        RECT 171.935 25.540 173.060 25.710 ;
        RECT 171.935 24.910 172.260 25.370 ;
        RECT 172.780 25.080 173.060 25.540 ;
        RECT 173.250 25.080 173.650 25.880 ;
        RECT 173.820 26.610 174.775 26.830 ;
        RECT 173.820 25.710 174.030 26.610 ;
        RECT 174.200 25.880 174.890 26.440 ;
        RECT 175.060 26.295 175.350 27.460 ;
        RECT 175.520 26.320 175.905 27.290 ;
        RECT 176.075 27.000 176.400 27.460 ;
        RECT 176.920 26.830 177.200 27.290 ;
        RECT 176.075 26.610 177.200 26.830 ;
        RECT 173.820 25.540 174.775 25.710 ;
        RECT 175.520 25.650 175.800 26.320 ;
        RECT 176.075 26.150 176.525 26.610 ;
        RECT 177.390 26.440 177.790 27.290 ;
        RECT 178.190 27.000 178.460 27.460 ;
        RECT 178.630 26.830 178.915 27.290 ;
        RECT 179.200 27.025 184.545 27.460 ;
        RECT 175.970 25.820 176.525 26.150 ;
        RECT 176.695 25.880 177.790 26.440 ;
        RECT 176.075 25.710 176.525 25.820 ;
        RECT 174.050 24.910 174.320 25.370 ;
        RECT 174.490 25.080 174.775 25.540 ;
        RECT 175.060 24.910 175.350 25.635 ;
        RECT 175.520 25.080 175.905 25.650 ;
        RECT 176.075 25.540 177.200 25.710 ;
        RECT 176.075 24.910 176.400 25.370 ;
        RECT 176.920 25.080 177.200 25.540 ;
        RECT 177.390 25.080 177.790 25.880 ;
        RECT 177.960 26.610 178.915 26.830 ;
        RECT 177.960 25.710 178.170 26.610 ;
        RECT 178.340 25.880 179.030 26.440 ;
        RECT 177.960 25.540 178.915 25.710 ;
        RECT 178.190 24.910 178.460 25.370 ;
        RECT 178.630 25.080 178.915 25.540 ;
        RECT 180.785 25.455 181.125 26.285 ;
        RECT 182.605 25.775 182.955 27.025 ;
        RECT 184.720 26.370 188.230 27.460 ;
        RECT 189.435 26.830 189.720 27.290 ;
        RECT 189.890 27.000 190.160 27.460 ;
        RECT 189.435 26.610 190.390 26.830 ;
        RECT 184.720 25.680 186.370 26.200 ;
        RECT 186.540 25.850 188.230 26.370 ;
        RECT 189.320 25.880 190.010 26.440 ;
        RECT 190.180 25.710 190.390 26.610 ;
        RECT 179.200 24.910 184.545 25.455 ;
        RECT 184.720 24.910 188.230 25.680 ;
        RECT 189.435 25.540 190.390 25.710 ;
        RECT 190.560 26.440 190.960 27.290 ;
        RECT 191.150 26.830 191.430 27.290 ;
        RECT 191.950 27.000 192.275 27.460 ;
        RECT 191.150 26.610 192.275 26.830 ;
        RECT 190.560 25.880 191.655 26.440 ;
        RECT 191.825 26.150 192.275 26.610 ;
        RECT 192.445 26.320 192.830 27.290 ;
        RECT 193.000 26.370 196.510 27.460 ;
        RECT 196.680 26.370 197.890 27.460 ;
        RECT 198.115 26.590 198.400 27.460 ;
        RECT 198.570 26.830 198.830 27.290 ;
        RECT 199.005 27.000 199.260 27.460 ;
        RECT 199.430 26.830 199.690 27.290 ;
        RECT 198.570 26.660 199.690 26.830 ;
        RECT 199.860 26.660 200.170 27.460 ;
        RECT 198.570 26.410 198.830 26.660 ;
        RECT 200.340 26.490 200.650 27.290 ;
        RECT 189.435 25.080 189.720 25.540 ;
        RECT 189.890 24.910 190.160 25.370 ;
        RECT 190.560 25.080 190.960 25.880 ;
        RECT 191.825 25.820 192.380 26.150 ;
        RECT 191.825 25.710 192.275 25.820 ;
        RECT 191.150 25.540 192.275 25.710 ;
        RECT 192.550 25.650 192.830 26.320 ;
        RECT 191.150 25.080 191.430 25.540 ;
        RECT 191.950 24.910 192.275 25.370 ;
        RECT 192.445 25.080 192.830 25.650 ;
        RECT 193.000 25.680 194.650 26.200 ;
        RECT 194.820 25.850 196.510 26.370 ;
        RECT 193.000 24.910 196.510 25.680 ;
        RECT 196.680 25.660 197.200 26.200 ;
        RECT 197.370 25.830 197.890 26.370 ;
        RECT 198.075 26.240 198.830 26.410 ;
        RECT 199.620 26.320 200.650 26.490 ;
        RECT 198.075 25.730 198.480 26.240 ;
        RECT 199.620 26.070 199.790 26.320 ;
        RECT 198.650 25.900 199.790 26.070 ;
        RECT 196.680 24.910 197.890 25.660 ;
        RECT 198.075 25.560 199.725 25.730 ;
        RECT 199.960 25.580 200.310 26.150 ;
        RECT 198.120 24.910 198.400 25.390 ;
        RECT 198.570 25.170 198.830 25.560 ;
        RECT 199.005 24.910 199.260 25.390 ;
        RECT 199.430 25.170 199.725 25.560 ;
        RECT 200.480 25.410 200.650 26.320 ;
        RECT 200.820 26.295 201.110 27.460 ;
        RECT 201.280 26.370 204.790 27.460 ;
        RECT 205.535 26.830 205.820 27.290 ;
        RECT 205.990 27.000 206.260 27.460 ;
        RECT 205.535 26.610 206.490 26.830 ;
        RECT 201.280 25.680 202.930 26.200 ;
        RECT 203.100 25.850 204.790 26.370 ;
        RECT 205.420 25.880 206.110 26.440 ;
        RECT 206.280 25.710 206.490 26.610 ;
        RECT 199.905 24.910 200.180 25.390 ;
        RECT 200.350 25.080 200.650 25.410 ;
        RECT 200.820 24.910 201.110 25.635 ;
        RECT 201.280 24.910 204.790 25.680 ;
        RECT 205.535 25.540 206.490 25.710 ;
        RECT 206.660 26.440 207.060 27.290 ;
        RECT 207.250 26.830 207.530 27.290 ;
        RECT 208.050 27.000 208.375 27.460 ;
        RECT 207.250 26.610 208.375 26.830 ;
        RECT 206.660 25.880 207.755 26.440 ;
        RECT 207.925 26.150 208.375 26.610 ;
        RECT 208.545 26.320 208.930 27.290 ;
        RECT 209.100 27.025 214.445 27.460 ;
        RECT 214.620 27.025 219.965 27.460 ;
        RECT 220.140 27.025 225.485 27.460 ;
        RECT 205.535 25.080 205.820 25.540 ;
        RECT 205.990 24.910 206.260 25.370 ;
        RECT 206.660 25.080 207.060 25.880 ;
        RECT 207.925 25.820 208.480 26.150 ;
        RECT 207.925 25.710 208.375 25.820 ;
        RECT 207.250 25.540 208.375 25.710 ;
        RECT 208.650 25.650 208.930 26.320 ;
        RECT 207.250 25.080 207.530 25.540 ;
        RECT 208.050 24.910 208.375 25.370 ;
        RECT 208.545 25.080 208.930 25.650 ;
        RECT 210.685 25.455 211.025 26.285 ;
        RECT 212.505 25.775 212.855 27.025 ;
        RECT 216.205 25.455 216.545 26.285 ;
        RECT 218.025 25.775 218.375 27.025 ;
        RECT 221.725 25.455 222.065 26.285 ;
        RECT 223.545 25.775 223.895 27.025 ;
        RECT 226.580 26.295 226.870 27.460 ;
        RECT 227.040 27.025 232.385 27.460 ;
        RECT 232.560 27.025 237.905 27.460 ;
        RECT 238.080 27.025 243.425 27.460 ;
        RECT 243.600 27.025 248.945 27.460 ;
        RECT 209.100 24.910 214.445 25.455 ;
        RECT 214.620 24.910 219.965 25.455 ;
        RECT 220.140 24.910 225.485 25.455 ;
        RECT 226.580 24.910 226.870 25.635 ;
        RECT 228.625 25.455 228.965 26.285 ;
        RECT 230.445 25.775 230.795 27.025 ;
        RECT 234.145 25.455 234.485 26.285 ;
        RECT 235.965 25.775 236.315 27.025 ;
        RECT 239.665 25.455 240.005 26.285 ;
        RECT 241.485 25.775 241.835 27.025 ;
        RECT 245.185 25.455 245.525 26.285 ;
        RECT 247.005 25.775 247.355 27.025 ;
        RECT 249.120 26.370 251.710 27.460 ;
        RECT 249.120 25.680 250.330 26.200 ;
        RECT 250.500 25.850 251.710 26.370 ;
        RECT 252.340 26.295 252.630 27.460 ;
        RECT 252.800 27.025 258.145 27.460 ;
        RECT 258.320 27.025 263.665 27.460 ;
        RECT 263.840 27.025 269.185 27.460 ;
        RECT 269.360 27.025 274.705 27.460 ;
        RECT 227.040 24.910 232.385 25.455 ;
        RECT 232.560 24.910 237.905 25.455 ;
        RECT 238.080 24.910 243.425 25.455 ;
        RECT 243.600 24.910 248.945 25.455 ;
        RECT 249.120 24.910 251.710 25.680 ;
        RECT 252.340 24.910 252.630 25.635 ;
        RECT 254.385 25.455 254.725 26.285 ;
        RECT 256.205 25.775 256.555 27.025 ;
        RECT 259.905 25.455 260.245 26.285 ;
        RECT 261.725 25.775 262.075 27.025 ;
        RECT 265.425 25.455 265.765 26.285 ;
        RECT 267.245 25.775 267.595 27.025 ;
        RECT 270.945 25.455 271.285 26.285 ;
        RECT 272.765 25.775 273.115 27.025 ;
        RECT 274.880 26.370 277.470 27.460 ;
        RECT 274.880 25.680 276.090 26.200 ;
        RECT 276.260 25.850 277.470 26.370 ;
        RECT 278.100 26.295 278.390 27.460 ;
        RECT 278.560 27.025 283.905 27.460 ;
        RECT 284.080 27.025 289.425 27.460 ;
        RECT 289.600 27.025 294.945 27.460 ;
        RECT 295.120 27.025 300.465 27.460 ;
        RECT 252.800 24.910 258.145 25.455 ;
        RECT 258.320 24.910 263.665 25.455 ;
        RECT 263.840 24.910 269.185 25.455 ;
        RECT 269.360 24.910 274.705 25.455 ;
        RECT 274.880 24.910 277.470 25.680 ;
        RECT 278.100 24.910 278.390 25.635 ;
        RECT 280.145 25.455 280.485 26.285 ;
        RECT 281.965 25.775 282.315 27.025 ;
        RECT 285.665 25.455 286.005 26.285 ;
        RECT 287.485 25.775 287.835 27.025 ;
        RECT 291.185 25.455 291.525 26.285 ;
        RECT 293.005 25.775 293.355 27.025 ;
        RECT 296.705 25.455 297.045 26.285 ;
        RECT 298.525 25.775 298.875 27.025 ;
        RECT 300.640 26.370 303.230 27.460 ;
        RECT 300.640 25.680 301.850 26.200 ;
        RECT 302.020 25.850 303.230 26.370 ;
        RECT 303.860 26.295 304.150 27.460 ;
        RECT 304.320 27.025 309.665 27.460 ;
        RECT 278.560 24.910 283.905 25.455 ;
        RECT 284.080 24.910 289.425 25.455 ;
        RECT 289.600 24.910 294.945 25.455 ;
        RECT 295.120 24.910 300.465 25.455 ;
        RECT 300.640 24.910 303.230 25.680 ;
        RECT 303.860 24.910 304.150 25.635 ;
        RECT 305.905 25.455 306.245 26.285 ;
        RECT 307.725 25.775 308.075 27.025 ;
        RECT 309.840 26.370 311.050 27.460 ;
        RECT 309.840 25.830 310.360 26.370 ;
        RECT 310.530 25.660 311.050 26.200 ;
        RECT 304.320 24.910 309.665 25.455 ;
        RECT 309.840 24.910 311.050 25.660 ;
        RECT 162.095 24.740 311.135 24.910 ;
        RECT 162.180 23.990 163.390 24.740 ;
        RECT 163.560 24.195 168.905 24.740 ;
        RECT 169.080 24.195 174.425 24.740 ;
        RECT 174.600 24.195 179.945 24.740 ;
        RECT 180.120 24.195 185.465 24.740 ;
        RECT 162.180 23.450 162.700 23.990 ;
        RECT 162.870 23.280 163.390 23.820 ;
        RECT 165.145 23.365 165.485 24.195 ;
        RECT 162.180 22.190 163.390 23.280 ;
        RECT 166.965 22.625 167.315 23.875 ;
        RECT 170.665 23.365 171.005 24.195 ;
        RECT 172.485 22.625 172.835 23.875 ;
        RECT 176.185 23.365 176.525 24.195 ;
        RECT 178.005 22.625 178.355 23.875 ;
        RECT 181.705 23.365 182.045 24.195 ;
        RECT 185.640 23.970 187.310 24.740 ;
        RECT 187.940 24.015 188.230 24.740 ;
        RECT 188.400 24.195 193.745 24.740 ;
        RECT 193.920 24.195 199.265 24.740 ;
        RECT 199.440 24.195 204.785 24.740 ;
        RECT 204.960 24.195 210.305 24.740 ;
        RECT 183.525 22.625 183.875 23.875 ;
        RECT 185.640 23.450 186.390 23.970 ;
        RECT 186.560 23.280 187.310 23.800 ;
        RECT 189.985 23.365 190.325 24.195 ;
        RECT 163.560 22.190 168.905 22.625 ;
        RECT 169.080 22.190 174.425 22.625 ;
        RECT 174.600 22.190 179.945 22.625 ;
        RECT 180.120 22.190 185.465 22.625 ;
        RECT 185.640 22.190 187.310 23.280 ;
        RECT 187.940 22.190 188.230 23.355 ;
        RECT 191.805 22.625 192.155 23.875 ;
        RECT 195.505 23.365 195.845 24.195 ;
        RECT 197.325 22.625 197.675 23.875 ;
        RECT 201.025 23.365 201.365 24.195 ;
        RECT 202.845 22.625 203.195 23.875 ;
        RECT 206.545 23.365 206.885 24.195 ;
        RECT 210.480 23.970 213.070 24.740 ;
        RECT 213.700 24.015 213.990 24.740 ;
        RECT 214.160 24.195 219.505 24.740 ;
        RECT 219.680 24.195 225.025 24.740 ;
        RECT 225.200 24.195 230.545 24.740 ;
        RECT 230.720 24.195 236.065 24.740 ;
        RECT 208.365 22.625 208.715 23.875 ;
        RECT 210.480 23.450 211.690 23.970 ;
        RECT 211.860 23.280 213.070 23.800 ;
        RECT 215.745 23.365 216.085 24.195 ;
        RECT 188.400 22.190 193.745 22.625 ;
        RECT 193.920 22.190 199.265 22.625 ;
        RECT 199.440 22.190 204.785 22.625 ;
        RECT 204.960 22.190 210.305 22.625 ;
        RECT 210.480 22.190 213.070 23.280 ;
        RECT 213.700 22.190 213.990 23.355 ;
        RECT 217.565 22.625 217.915 23.875 ;
        RECT 221.265 23.365 221.605 24.195 ;
        RECT 223.085 22.625 223.435 23.875 ;
        RECT 226.785 23.365 227.125 24.195 ;
        RECT 228.605 22.625 228.955 23.875 ;
        RECT 232.305 23.365 232.645 24.195 ;
        RECT 236.240 23.970 238.830 24.740 ;
        RECT 239.460 24.015 239.750 24.740 ;
        RECT 239.920 24.195 245.265 24.740 ;
        RECT 245.440 24.195 250.785 24.740 ;
        RECT 250.960 24.195 256.305 24.740 ;
        RECT 256.480 24.195 261.825 24.740 ;
        RECT 234.125 22.625 234.475 23.875 ;
        RECT 236.240 23.450 237.450 23.970 ;
        RECT 237.620 23.280 238.830 23.800 ;
        RECT 241.505 23.365 241.845 24.195 ;
        RECT 214.160 22.190 219.505 22.625 ;
        RECT 219.680 22.190 225.025 22.625 ;
        RECT 225.200 22.190 230.545 22.625 ;
        RECT 230.720 22.190 236.065 22.625 ;
        RECT 236.240 22.190 238.830 23.280 ;
        RECT 239.460 22.190 239.750 23.355 ;
        RECT 243.325 22.625 243.675 23.875 ;
        RECT 247.025 23.365 247.365 24.195 ;
        RECT 248.845 22.625 249.195 23.875 ;
        RECT 252.545 23.365 252.885 24.195 ;
        RECT 254.365 22.625 254.715 23.875 ;
        RECT 258.065 23.365 258.405 24.195 ;
        RECT 262.000 23.970 264.590 24.740 ;
        RECT 265.220 24.015 265.510 24.740 ;
        RECT 265.680 24.195 271.025 24.740 ;
        RECT 271.200 24.195 276.545 24.740 ;
        RECT 276.720 24.195 282.065 24.740 ;
        RECT 282.240 24.195 287.585 24.740 ;
        RECT 259.885 22.625 260.235 23.875 ;
        RECT 262.000 23.450 263.210 23.970 ;
        RECT 263.380 23.280 264.590 23.800 ;
        RECT 267.265 23.365 267.605 24.195 ;
        RECT 239.920 22.190 245.265 22.625 ;
        RECT 245.440 22.190 250.785 22.625 ;
        RECT 250.960 22.190 256.305 22.625 ;
        RECT 256.480 22.190 261.825 22.625 ;
        RECT 262.000 22.190 264.590 23.280 ;
        RECT 265.220 22.190 265.510 23.355 ;
        RECT 269.085 22.625 269.435 23.875 ;
        RECT 272.785 23.365 273.125 24.195 ;
        RECT 274.605 22.625 274.955 23.875 ;
        RECT 278.305 23.365 278.645 24.195 ;
        RECT 280.125 22.625 280.475 23.875 ;
        RECT 283.825 23.365 284.165 24.195 ;
        RECT 287.760 23.970 290.350 24.740 ;
        RECT 290.980 24.015 291.270 24.740 ;
        RECT 291.440 24.195 296.785 24.740 ;
        RECT 296.960 24.195 302.305 24.740 ;
        RECT 302.480 24.195 307.825 24.740 ;
        RECT 285.645 22.625 285.995 23.875 ;
        RECT 287.760 23.450 288.970 23.970 ;
        RECT 289.140 23.280 290.350 23.800 ;
        RECT 293.025 23.365 293.365 24.195 ;
        RECT 265.680 22.190 271.025 22.625 ;
        RECT 271.200 22.190 276.545 22.625 ;
        RECT 276.720 22.190 282.065 22.625 ;
        RECT 282.240 22.190 287.585 22.625 ;
        RECT 287.760 22.190 290.350 23.280 ;
        RECT 290.980 22.190 291.270 23.355 ;
        RECT 294.845 22.625 295.195 23.875 ;
        RECT 298.545 23.365 298.885 24.195 ;
        RECT 300.365 22.625 300.715 23.875 ;
        RECT 304.065 23.365 304.405 24.195 ;
        RECT 308.000 23.970 309.670 24.740 ;
        RECT 309.840 23.990 311.050 24.740 ;
        RECT 305.885 22.625 306.235 23.875 ;
        RECT 308.000 23.450 308.750 23.970 ;
        RECT 308.920 23.280 309.670 23.800 ;
        RECT 291.440 22.190 296.785 22.625 ;
        RECT 296.960 22.190 302.305 22.625 ;
        RECT 302.480 22.190 307.825 22.625 ;
        RECT 308.000 22.190 309.670 23.280 ;
        RECT 309.840 23.280 310.360 23.820 ;
        RECT 310.530 23.450 311.050 23.990 ;
        RECT 309.840 22.190 311.050 23.280 ;
        RECT 162.095 22.020 311.135 22.190 ;
        RECT 162.180 20.930 163.390 22.020 ;
        RECT 163.560 21.585 168.905 22.020 ;
        RECT 169.080 21.585 174.425 22.020 ;
        RECT 162.180 20.220 162.700 20.760 ;
        RECT 162.870 20.390 163.390 20.930 ;
        RECT 162.180 19.470 163.390 20.220 ;
        RECT 165.145 20.015 165.485 20.845 ;
        RECT 166.965 20.335 167.315 21.585 ;
        RECT 170.665 20.015 171.005 20.845 ;
        RECT 172.485 20.335 172.835 21.585 ;
        RECT 175.060 20.855 175.350 22.020 ;
        RECT 175.520 21.585 180.865 22.020 ;
        RECT 181.040 21.585 186.385 22.020 ;
        RECT 186.560 21.585 191.905 22.020 ;
        RECT 192.080 21.585 197.425 22.020 ;
        RECT 163.560 19.470 168.905 20.015 ;
        RECT 169.080 19.470 174.425 20.015 ;
        RECT 175.060 19.470 175.350 20.195 ;
        RECT 177.105 20.015 177.445 20.845 ;
        RECT 178.925 20.335 179.275 21.585 ;
        RECT 182.625 20.015 182.965 20.845 ;
        RECT 184.445 20.335 184.795 21.585 ;
        RECT 188.145 20.015 188.485 20.845 ;
        RECT 189.965 20.335 190.315 21.585 ;
        RECT 193.665 20.015 194.005 20.845 ;
        RECT 195.485 20.335 195.835 21.585 ;
        RECT 197.600 20.930 200.190 22.020 ;
        RECT 197.600 20.240 198.810 20.760 ;
        RECT 198.980 20.410 200.190 20.930 ;
        RECT 200.820 20.855 201.110 22.020 ;
        RECT 201.280 21.585 206.625 22.020 ;
        RECT 206.800 21.585 212.145 22.020 ;
        RECT 212.320 21.585 217.665 22.020 ;
        RECT 217.840 21.585 223.185 22.020 ;
        RECT 175.520 19.470 180.865 20.015 ;
        RECT 181.040 19.470 186.385 20.015 ;
        RECT 186.560 19.470 191.905 20.015 ;
        RECT 192.080 19.470 197.425 20.015 ;
        RECT 197.600 19.470 200.190 20.240 ;
        RECT 200.820 19.470 201.110 20.195 ;
        RECT 202.865 20.015 203.205 20.845 ;
        RECT 204.685 20.335 205.035 21.585 ;
        RECT 208.385 20.015 208.725 20.845 ;
        RECT 210.205 20.335 210.555 21.585 ;
        RECT 213.905 20.015 214.245 20.845 ;
        RECT 215.725 20.335 216.075 21.585 ;
        RECT 219.425 20.015 219.765 20.845 ;
        RECT 221.245 20.335 221.595 21.585 ;
        RECT 223.360 20.930 225.950 22.020 ;
        RECT 223.360 20.240 224.570 20.760 ;
        RECT 224.740 20.410 225.950 20.930 ;
        RECT 226.580 20.855 226.870 22.020 ;
        RECT 227.040 21.585 232.385 22.020 ;
        RECT 232.560 21.585 237.905 22.020 ;
        RECT 238.080 21.585 243.425 22.020 ;
        RECT 243.600 21.585 248.945 22.020 ;
        RECT 201.280 19.470 206.625 20.015 ;
        RECT 206.800 19.470 212.145 20.015 ;
        RECT 212.320 19.470 217.665 20.015 ;
        RECT 217.840 19.470 223.185 20.015 ;
        RECT 223.360 19.470 225.950 20.240 ;
        RECT 226.580 19.470 226.870 20.195 ;
        RECT 228.625 20.015 228.965 20.845 ;
        RECT 230.445 20.335 230.795 21.585 ;
        RECT 234.145 20.015 234.485 20.845 ;
        RECT 235.965 20.335 236.315 21.585 ;
        RECT 239.665 20.015 240.005 20.845 ;
        RECT 241.485 20.335 241.835 21.585 ;
        RECT 245.185 20.015 245.525 20.845 ;
        RECT 247.005 20.335 247.355 21.585 ;
        RECT 249.120 20.930 251.710 22.020 ;
        RECT 249.120 20.240 250.330 20.760 ;
        RECT 250.500 20.410 251.710 20.930 ;
        RECT 252.340 20.855 252.630 22.020 ;
        RECT 252.800 21.585 258.145 22.020 ;
        RECT 258.320 21.585 263.665 22.020 ;
        RECT 263.840 21.585 269.185 22.020 ;
        RECT 269.360 21.585 274.705 22.020 ;
        RECT 227.040 19.470 232.385 20.015 ;
        RECT 232.560 19.470 237.905 20.015 ;
        RECT 238.080 19.470 243.425 20.015 ;
        RECT 243.600 19.470 248.945 20.015 ;
        RECT 249.120 19.470 251.710 20.240 ;
        RECT 252.340 19.470 252.630 20.195 ;
        RECT 254.385 20.015 254.725 20.845 ;
        RECT 256.205 20.335 256.555 21.585 ;
        RECT 259.905 20.015 260.245 20.845 ;
        RECT 261.725 20.335 262.075 21.585 ;
        RECT 265.425 20.015 265.765 20.845 ;
        RECT 267.245 20.335 267.595 21.585 ;
        RECT 270.945 20.015 271.285 20.845 ;
        RECT 272.765 20.335 273.115 21.585 ;
        RECT 274.880 20.930 277.470 22.020 ;
        RECT 274.880 20.240 276.090 20.760 ;
        RECT 276.260 20.410 277.470 20.930 ;
        RECT 278.100 20.855 278.390 22.020 ;
        RECT 278.560 21.585 283.905 22.020 ;
        RECT 284.080 21.585 289.425 22.020 ;
        RECT 289.600 21.585 294.945 22.020 ;
        RECT 295.120 21.585 300.465 22.020 ;
        RECT 252.800 19.470 258.145 20.015 ;
        RECT 258.320 19.470 263.665 20.015 ;
        RECT 263.840 19.470 269.185 20.015 ;
        RECT 269.360 19.470 274.705 20.015 ;
        RECT 274.880 19.470 277.470 20.240 ;
        RECT 278.100 19.470 278.390 20.195 ;
        RECT 280.145 20.015 280.485 20.845 ;
        RECT 281.965 20.335 282.315 21.585 ;
        RECT 285.665 20.015 286.005 20.845 ;
        RECT 287.485 20.335 287.835 21.585 ;
        RECT 291.185 20.015 291.525 20.845 ;
        RECT 293.005 20.335 293.355 21.585 ;
        RECT 296.705 20.015 297.045 20.845 ;
        RECT 298.525 20.335 298.875 21.585 ;
        RECT 300.640 20.930 303.230 22.020 ;
        RECT 300.640 20.240 301.850 20.760 ;
        RECT 302.020 20.410 303.230 20.930 ;
        RECT 303.860 20.855 304.150 22.020 ;
        RECT 304.320 21.585 309.665 22.020 ;
        RECT 278.560 19.470 283.905 20.015 ;
        RECT 284.080 19.470 289.425 20.015 ;
        RECT 289.600 19.470 294.945 20.015 ;
        RECT 295.120 19.470 300.465 20.015 ;
        RECT 300.640 19.470 303.230 20.240 ;
        RECT 303.860 19.470 304.150 20.195 ;
        RECT 305.905 20.015 306.245 20.845 ;
        RECT 307.725 20.335 308.075 21.585 ;
        RECT 309.840 20.930 311.050 22.020 ;
        RECT 309.840 20.390 310.360 20.930 ;
        RECT 310.530 20.220 311.050 20.760 ;
        RECT 304.320 19.470 309.665 20.015 ;
        RECT 309.840 19.470 311.050 20.220 ;
        RECT 162.095 19.300 311.135 19.470 ;
        RECT 162.180 18.550 163.390 19.300 ;
        RECT 163.560 18.755 168.905 19.300 ;
        RECT 169.080 18.755 174.425 19.300 ;
        RECT 174.600 18.755 179.945 19.300 ;
        RECT 180.120 18.755 185.465 19.300 ;
        RECT 162.180 18.010 162.700 18.550 ;
        RECT 162.870 17.840 163.390 18.380 ;
        RECT 165.145 17.925 165.485 18.755 ;
        RECT 162.180 16.750 163.390 17.840 ;
        RECT 166.965 17.185 167.315 18.435 ;
        RECT 170.665 17.925 171.005 18.755 ;
        RECT 172.485 17.185 172.835 18.435 ;
        RECT 176.185 17.925 176.525 18.755 ;
        RECT 178.005 17.185 178.355 18.435 ;
        RECT 181.705 17.925 182.045 18.755 ;
        RECT 185.640 18.530 187.310 19.300 ;
        RECT 187.940 18.575 188.230 19.300 ;
        RECT 188.400 18.755 193.745 19.300 ;
        RECT 193.920 18.755 199.265 19.300 ;
        RECT 199.440 18.755 204.785 19.300 ;
        RECT 204.960 18.755 210.305 19.300 ;
        RECT 183.525 17.185 183.875 18.435 ;
        RECT 185.640 18.010 186.390 18.530 ;
        RECT 186.560 17.840 187.310 18.360 ;
        RECT 189.985 17.925 190.325 18.755 ;
        RECT 163.560 16.750 168.905 17.185 ;
        RECT 169.080 16.750 174.425 17.185 ;
        RECT 174.600 16.750 179.945 17.185 ;
        RECT 180.120 16.750 185.465 17.185 ;
        RECT 185.640 16.750 187.310 17.840 ;
        RECT 187.940 16.750 188.230 17.915 ;
        RECT 191.805 17.185 192.155 18.435 ;
        RECT 195.505 17.925 195.845 18.755 ;
        RECT 197.325 17.185 197.675 18.435 ;
        RECT 201.025 17.925 201.365 18.755 ;
        RECT 202.845 17.185 203.195 18.435 ;
        RECT 206.545 17.925 206.885 18.755 ;
        RECT 210.480 18.530 213.070 19.300 ;
        RECT 213.700 18.575 213.990 19.300 ;
        RECT 214.160 18.755 219.505 19.300 ;
        RECT 219.680 18.755 225.025 19.300 ;
        RECT 225.200 18.755 230.545 19.300 ;
        RECT 230.720 18.755 236.065 19.300 ;
        RECT 208.365 17.185 208.715 18.435 ;
        RECT 210.480 18.010 211.690 18.530 ;
        RECT 211.860 17.840 213.070 18.360 ;
        RECT 215.745 17.925 216.085 18.755 ;
        RECT 188.400 16.750 193.745 17.185 ;
        RECT 193.920 16.750 199.265 17.185 ;
        RECT 199.440 16.750 204.785 17.185 ;
        RECT 204.960 16.750 210.305 17.185 ;
        RECT 210.480 16.750 213.070 17.840 ;
        RECT 213.700 16.750 213.990 17.915 ;
        RECT 217.565 17.185 217.915 18.435 ;
        RECT 221.265 17.925 221.605 18.755 ;
        RECT 223.085 17.185 223.435 18.435 ;
        RECT 226.785 17.925 227.125 18.755 ;
        RECT 228.605 17.185 228.955 18.435 ;
        RECT 232.305 17.925 232.645 18.755 ;
        RECT 236.240 18.530 238.830 19.300 ;
        RECT 239.460 18.575 239.750 19.300 ;
        RECT 239.920 18.755 245.265 19.300 ;
        RECT 245.440 18.755 250.785 19.300 ;
        RECT 250.960 18.755 256.305 19.300 ;
        RECT 256.480 18.755 261.825 19.300 ;
        RECT 234.125 17.185 234.475 18.435 ;
        RECT 236.240 18.010 237.450 18.530 ;
        RECT 237.620 17.840 238.830 18.360 ;
        RECT 241.505 17.925 241.845 18.755 ;
        RECT 214.160 16.750 219.505 17.185 ;
        RECT 219.680 16.750 225.025 17.185 ;
        RECT 225.200 16.750 230.545 17.185 ;
        RECT 230.720 16.750 236.065 17.185 ;
        RECT 236.240 16.750 238.830 17.840 ;
        RECT 239.460 16.750 239.750 17.915 ;
        RECT 243.325 17.185 243.675 18.435 ;
        RECT 247.025 17.925 247.365 18.755 ;
        RECT 248.845 17.185 249.195 18.435 ;
        RECT 252.545 17.925 252.885 18.755 ;
        RECT 254.365 17.185 254.715 18.435 ;
        RECT 258.065 17.925 258.405 18.755 ;
        RECT 262.000 18.530 264.590 19.300 ;
        RECT 265.220 18.575 265.510 19.300 ;
        RECT 265.680 18.755 271.025 19.300 ;
        RECT 271.200 18.755 276.545 19.300 ;
        RECT 276.720 18.755 282.065 19.300 ;
        RECT 282.240 18.755 287.585 19.300 ;
        RECT 259.885 17.185 260.235 18.435 ;
        RECT 262.000 18.010 263.210 18.530 ;
        RECT 263.380 17.840 264.590 18.360 ;
        RECT 267.265 17.925 267.605 18.755 ;
        RECT 239.920 16.750 245.265 17.185 ;
        RECT 245.440 16.750 250.785 17.185 ;
        RECT 250.960 16.750 256.305 17.185 ;
        RECT 256.480 16.750 261.825 17.185 ;
        RECT 262.000 16.750 264.590 17.840 ;
        RECT 265.220 16.750 265.510 17.915 ;
        RECT 269.085 17.185 269.435 18.435 ;
        RECT 272.785 17.925 273.125 18.755 ;
        RECT 274.605 17.185 274.955 18.435 ;
        RECT 278.305 17.925 278.645 18.755 ;
        RECT 280.125 17.185 280.475 18.435 ;
        RECT 283.825 17.925 284.165 18.755 ;
        RECT 287.760 18.530 290.350 19.300 ;
        RECT 290.980 18.575 291.270 19.300 ;
        RECT 291.440 18.755 296.785 19.300 ;
        RECT 296.960 18.755 302.305 19.300 ;
        RECT 302.480 18.755 307.825 19.300 ;
        RECT 285.645 17.185 285.995 18.435 ;
        RECT 287.760 18.010 288.970 18.530 ;
        RECT 289.140 17.840 290.350 18.360 ;
        RECT 293.025 17.925 293.365 18.755 ;
        RECT 265.680 16.750 271.025 17.185 ;
        RECT 271.200 16.750 276.545 17.185 ;
        RECT 276.720 16.750 282.065 17.185 ;
        RECT 282.240 16.750 287.585 17.185 ;
        RECT 287.760 16.750 290.350 17.840 ;
        RECT 290.980 16.750 291.270 17.915 ;
        RECT 294.845 17.185 295.195 18.435 ;
        RECT 298.545 17.925 298.885 18.755 ;
        RECT 300.365 17.185 300.715 18.435 ;
        RECT 304.065 17.925 304.405 18.755 ;
        RECT 308.000 18.530 309.670 19.300 ;
        RECT 309.840 18.550 311.050 19.300 ;
        RECT 305.885 17.185 306.235 18.435 ;
        RECT 308.000 18.010 308.750 18.530 ;
        RECT 308.920 17.840 309.670 18.360 ;
        RECT 291.440 16.750 296.785 17.185 ;
        RECT 296.960 16.750 302.305 17.185 ;
        RECT 302.480 16.750 307.825 17.185 ;
        RECT 308.000 16.750 309.670 17.840 ;
        RECT 309.840 17.840 310.360 18.380 ;
        RECT 310.530 18.010 311.050 18.550 ;
        RECT 309.840 16.750 311.050 17.840 ;
        RECT 162.095 16.580 311.135 16.750 ;
        RECT 162.180 15.490 163.390 16.580 ;
        RECT 163.560 16.145 168.905 16.580 ;
        RECT 169.080 16.145 174.425 16.580 ;
        RECT 162.180 14.780 162.700 15.320 ;
        RECT 162.870 14.950 163.390 15.490 ;
        RECT 162.180 14.030 163.390 14.780 ;
        RECT 165.145 14.575 165.485 15.405 ;
        RECT 166.965 14.895 167.315 16.145 ;
        RECT 170.665 14.575 171.005 15.405 ;
        RECT 172.485 14.895 172.835 16.145 ;
        RECT 175.060 15.415 175.350 16.580 ;
        RECT 175.520 16.145 180.865 16.580 ;
        RECT 181.040 16.145 186.385 16.580 ;
        RECT 163.560 14.030 168.905 14.575 ;
        RECT 169.080 14.030 174.425 14.575 ;
        RECT 175.060 14.030 175.350 14.755 ;
        RECT 177.105 14.575 177.445 15.405 ;
        RECT 178.925 14.895 179.275 16.145 ;
        RECT 182.625 14.575 182.965 15.405 ;
        RECT 184.445 14.895 184.795 16.145 ;
        RECT 186.560 15.490 187.770 16.580 ;
        RECT 186.560 14.780 187.080 15.320 ;
        RECT 187.250 14.950 187.770 15.490 ;
        RECT 187.940 15.415 188.230 16.580 ;
        RECT 188.400 16.145 193.745 16.580 ;
        RECT 193.920 16.145 199.265 16.580 ;
        RECT 175.520 14.030 180.865 14.575 ;
        RECT 181.040 14.030 186.385 14.575 ;
        RECT 186.560 14.030 187.770 14.780 ;
        RECT 187.940 14.030 188.230 14.755 ;
        RECT 189.985 14.575 190.325 15.405 ;
        RECT 191.805 14.895 192.155 16.145 ;
        RECT 195.505 14.575 195.845 15.405 ;
        RECT 197.325 14.895 197.675 16.145 ;
        RECT 199.440 15.490 200.650 16.580 ;
        RECT 199.440 14.780 199.960 15.320 ;
        RECT 200.130 14.950 200.650 15.490 ;
        RECT 200.820 15.415 201.110 16.580 ;
        RECT 201.280 16.145 206.625 16.580 ;
        RECT 206.800 16.145 212.145 16.580 ;
        RECT 188.400 14.030 193.745 14.575 ;
        RECT 193.920 14.030 199.265 14.575 ;
        RECT 199.440 14.030 200.650 14.780 ;
        RECT 200.820 14.030 201.110 14.755 ;
        RECT 202.865 14.575 203.205 15.405 ;
        RECT 204.685 14.895 205.035 16.145 ;
        RECT 208.385 14.575 208.725 15.405 ;
        RECT 210.205 14.895 210.555 16.145 ;
        RECT 212.320 15.490 213.530 16.580 ;
        RECT 212.320 14.780 212.840 15.320 ;
        RECT 213.010 14.950 213.530 15.490 ;
        RECT 213.700 15.415 213.990 16.580 ;
        RECT 214.160 16.145 219.505 16.580 ;
        RECT 219.680 16.145 225.025 16.580 ;
        RECT 201.280 14.030 206.625 14.575 ;
        RECT 206.800 14.030 212.145 14.575 ;
        RECT 212.320 14.030 213.530 14.780 ;
        RECT 213.700 14.030 213.990 14.755 ;
        RECT 215.745 14.575 216.085 15.405 ;
        RECT 217.565 14.895 217.915 16.145 ;
        RECT 221.265 14.575 221.605 15.405 ;
        RECT 223.085 14.895 223.435 16.145 ;
        RECT 225.200 15.490 226.410 16.580 ;
        RECT 225.200 14.780 225.720 15.320 ;
        RECT 225.890 14.950 226.410 15.490 ;
        RECT 226.580 15.415 226.870 16.580 ;
        RECT 227.040 16.145 232.385 16.580 ;
        RECT 232.560 16.145 237.905 16.580 ;
        RECT 214.160 14.030 219.505 14.575 ;
        RECT 219.680 14.030 225.025 14.575 ;
        RECT 225.200 14.030 226.410 14.780 ;
        RECT 226.580 14.030 226.870 14.755 ;
        RECT 228.625 14.575 228.965 15.405 ;
        RECT 230.445 14.895 230.795 16.145 ;
        RECT 234.145 14.575 234.485 15.405 ;
        RECT 235.965 14.895 236.315 16.145 ;
        RECT 238.080 15.490 239.290 16.580 ;
        RECT 238.080 14.780 238.600 15.320 ;
        RECT 238.770 14.950 239.290 15.490 ;
        RECT 239.460 15.415 239.750 16.580 ;
        RECT 239.920 16.145 245.265 16.580 ;
        RECT 245.440 16.145 250.785 16.580 ;
        RECT 227.040 14.030 232.385 14.575 ;
        RECT 232.560 14.030 237.905 14.575 ;
        RECT 238.080 14.030 239.290 14.780 ;
        RECT 239.460 14.030 239.750 14.755 ;
        RECT 241.505 14.575 241.845 15.405 ;
        RECT 243.325 14.895 243.675 16.145 ;
        RECT 247.025 14.575 247.365 15.405 ;
        RECT 248.845 14.895 249.195 16.145 ;
        RECT 250.960 15.490 252.170 16.580 ;
        RECT 250.960 14.780 251.480 15.320 ;
        RECT 251.650 14.950 252.170 15.490 ;
        RECT 252.340 15.415 252.630 16.580 ;
        RECT 252.800 16.145 258.145 16.580 ;
        RECT 258.320 16.145 263.665 16.580 ;
        RECT 239.920 14.030 245.265 14.575 ;
        RECT 245.440 14.030 250.785 14.575 ;
        RECT 250.960 14.030 252.170 14.780 ;
        RECT 252.340 14.030 252.630 14.755 ;
        RECT 254.385 14.575 254.725 15.405 ;
        RECT 256.205 14.895 256.555 16.145 ;
        RECT 259.905 14.575 260.245 15.405 ;
        RECT 261.725 14.895 262.075 16.145 ;
        RECT 263.840 15.490 265.050 16.580 ;
        RECT 263.840 14.780 264.360 15.320 ;
        RECT 264.530 14.950 265.050 15.490 ;
        RECT 265.220 15.415 265.510 16.580 ;
        RECT 265.680 16.145 271.025 16.580 ;
        RECT 271.200 16.145 276.545 16.580 ;
        RECT 252.800 14.030 258.145 14.575 ;
        RECT 258.320 14.030 263.665 14.575 ;
        RECT 263.840 14.030 265.050 14.780 ;
        RECT 265.220 14.030 265.510 14.755 ;
        RECT 267.265 14.575 267.605 15.405 ;
        RECT 269.085 14.895 269.435 16.145 ;
        RECT 272.785 14.575 273.125 15.405 ;
        RECT 274.605 14.895 274.955 16.145 ;
        RECT 276.720 15.490 277.930 16.580 ;
        RECT 276.720 14.780 277.240 15.320 ;
        RECT 277.410 14.950 277.930 15.490 ;
        RECT 278.100 15.415 278.390 16.580 ;
        RECT 278.560 16.145 283.905 16.580 ;
        RECT 284.080 16.145 289.425 16.580 ;
        RECT 265.680 14.030 271.025 14.575 ;
        RECT 271.200 14.030 276.545 14.575 ;
        RECT 276.720 14.030 277.930 14.780 ;
        RECT 278.100 14.030 278.390 14.755 ;
        RECT 280.145 14.575 280.485 15.405 ;
        RECT 281.965 14.895 282.315 16.145 ;
        RECT 285.665 14.575 286.005 15.405 ;
        RECT 287.485 14.895 287.835 16.145 ;
        RECT 289.600 15.490 290.810 16.580 ;
        RECT 289.600 14.780 290.120 15.320 ;
        RECT 290.290 14.950 290.810 15.490 ;
        RECT 290.980 15.415 291.270 16.580 ;
        RECT 291.440 16.145 296.785 16.580 ;
        RECT 296.960 16.145 302.305 16.580 ;
        RECT 278.560 14.030 283.905 14.575 ;
        RECT 284.080 14.030 289.425 14.575 ;
        RECT 289.600 14.030 290.810 14.780 ;
        RECT 290.980 14.030 291.270 14.755 ;
        RECT 293.025 14.575 293.365 15.405 ;
        RECT 294.845 14.895 295.195 16.145 ;
        RECT 298.545 14.575 298.885 15.405 ;
        RECT 300.365 14.895 300.715 16.145 ;
        RECT 302.480 15.490 303.690 16.580 ;
        RECT 302.480 14.780 303.000 15.320 ;
        RECT 303.170 14.950 303.690 15.490 ;
        RECT 303.860 15.415 304.150 16.580 ;
        RECT 304.320 16.145 309.665 16.580 ;
        RECT 291.440 14.030 296.785 14.575 ;
        RECT 296.960 14.030 302.305 14.575 ;
        RECT 302.480 14.030 303.690 14.780 ;
        RECT 303.860 14.030 304.150 14.755 ;
        RECT 305.905 14.575 306.245 15.405 ;
        RECT 307.725 14.895 308.075 16.145 ;
        RECT 309.840 15.490 311.050 16.580 ;
        RECT 309.840 14.950 310.360 15.490 ;
        RECT 310.530 14.780 311.050 15.320 ;
        RECT 304.320 14.030 309.665 14.575 ;
        RECT 309.840 14.030 311.050 14.780 ;
        RECT 162.095 13.860 311.135 14.030 ;
        RECT 4.300 4.300 155.700 4.700 ;
      LAYER met1 ;
        RECT 45.390 225.410 246.965 225.710 ;
        RECT 45.390 224.810 45.690 225.410 ;
        RECT 59.190 224.810 236.370 225.110 ;
        RECT 246.665 225.010 246.965 225.410 ;
        RECT 62.000 224.210 226.710 224.510 ;
        RECT 236.070 224.410 236.370 224.810 ;
        RECT 226.410 223.810 226.710 224.210 ;
        RECT 4.100 216.515 102.825 222.630 ;
        RECT 106.340 220.315 153.245 220.715 ;
        RECT 106.340 217.515 108.920 220.315 ;
        RECT 109.605 219.705 110.565 219.935 ;
        RECT 110.895 219.705 111.855 220.055 ;
        RECT 109.325 219.255 109.555 219.500 ;
        RECT 110.615 219.255 110.845 219.500 ;
        RECT 111.905 219.255 112.135 219.500 ;
        RECT 109.290 217.755 109.590 219.255 ;
        RECT 110.580 217.755 110.880 219.255 ;
        RECT 111.870 217.755 112.170 219.255 ;
        RECT 4.100 212.490 63.455 216.515 ;
        RECT 64.175 215.825 80.135 216.055 ;
        RECT 81.805 215.825 97.765 216.055 ;
        RECT 63.895 214.620 64.125 215.620 ;
        RECT 80.185 214.620 81.755 215.620 ;
        RECT 97.815 214.620 98.045 215.620 ;
        RECT 64.175 214.185 80.135 214.415 ;
        RECT 81.805 214.185 97.765 214.415 ;
        RECT 77.595 213.035 78.595 213.270 ;
        RECT 83.345 213.035 84.345 213.270 ;
        RECT 64.175 212.805 80.135 213.035 ;
        RECT 81.805 212.805 97.765 213.035 ;
        RECT 4.100 211.660 56.570 212.490 ;
        RECT 4.100 191.850 9.525 211.660 ;
        RECT 10.245 210.970 18.205 211.200 ;
        RECT 18.535 210.970 26.495 211.200 ;
        RECT 28.165 210.970 36.125 211.200 ;
        RECT 36.455 210.970 44.415 211.200 ;
        RECT 9.965 210.465 10.195 210.765 ;
        RECT 9.925 209.065 10.225 210.465 ;
        RECT 9.965 202.765 10.195 209.065 ;
        RECT 18.255 207.465 18.485 210.765 ;
        RECT 18.215 206.065 18.515 207.465 ;
        RECT 18.255 202.765 18.485 206.065 ;
        RECT 26.545 204.465 26.775 210.765 ;
        RECT 27.885 204.465 28.115 210.765 ;
        RECT 36.175 207.465 36.405 210.765 ;
        RECT 44.465 210.465 44.695 210.765 ;
        RECT 44.425 209.065 44.725 210.465 ;
        RECT 45.135 210.150 56.570 211.660 ;
        RECT 36.165 206.065 36.465 207.465 ;
        RECT 26.505 203.065 26.805 204.465 ;
        RECT 27.845 203.065 28.145 204.465 ;
        RECT 26.505 202.560 28.145 203.065 ;
        RECT 36.175 202.765 36.405 206.065 ;
        RECT 44.465 202.765 44.695 209.065 ;
        RECT 45.135 207.460 50.745 210.150 ;
        RECT 54.835 209.565 56.570 210.150 ;
        RECT 51.315 207.460 51.905 209.565 ;
        RECT 52.485 207.460 54.245 209.565 ;
        RECT 54.825 207.460 56.570 209.565 ;
        RECT 10.245 202.330 18.205 202.560 ;
        RECT 18.535 202.330 36.125 202.560 ;
        RECT 36.455 202.330 44.415 202.560 ;
        RECT 10.245 201.180 44.415 202.330 ;
        RECT 10.245 200.950 18.205 201.180 ;
        RECT 18.535 200.950 36.125 201.180 ;
        RECT 36.455 200.950 44.415 201.180 ;
        RECT 9.965 194.445 10.195 200.745 ;
        RECT 18.255 197.445 18.485 200.745 ;
        RECT 26.505 200.445 28.145 200.950 ;
        RECT 26.505 199.045 26.805 200.445 ;
        RECT 27.845 199.045 28.145 200.445 ;
        RECT 18.215 196.045 18.515 197.445 ;
        RECT 9.925 193.045 10.225 194.445 ;
        RECT 9.965 192.745 10.195 193.045 ;
        RECT 18.255 192.745 18.485 196.045 ;
        RECT 26.545 192.745 26.775 199.045 ;
        RECT 27.885 192.745 28.115 199.045 ;
        RECT 36.175 197.445 36.405 200.745 ;
        RECT 36.165 196.045 36.465 197.445 ;
        RECT 36.175 192.745 36.405 196.045 ;
        RECT 44.465 194.445 44.695 200.745 ;
        RECT 44.425 193.045 44.725 194.445 ;
        RECT 44.465 192.745 44.695 193.045 ;
        RECT 10.245 192.310 18.205 192.540 ;
        RECT 18.535 192.310 26.495 192.540 ;
        RECT 28.165 192.310 36.125 192.540 ;
        RECT 36.455 192.310 44.415 192.540 ;
        RECT 45.135 191.850 49.450 207.460 ;
        RECT 4.100 190.670 49.450 191.850 ;
        RECT 4.100 180.880 9.525 190.670 ;
        RECT 9.965 189.980 12.205 190.210 ;
        RECT 12.535 189.980 14.495 190.210 ;
        RECT 9.965 184.050 10.195 189.980 ;
        RECT 12.535 189.775 13.090 189.980 ;
        RECT 12.255 189.350 13.090 189.775 ;
        RECT 9.930 182.650 10.230 184.050 ;
        RECT 9.965 181.570 10.195 182.650 ;
        RECT 12.255 181.775 12.485 189.350 ;
        RECT 14.545 188.900 14.775 189.775 ;
        RECT 14.510 187.500 14.810 188.900 ;
        RECT 14.545 181.775 14.775 187.500 ;
        RECT 9.965 181.340 12.205 181.570 ;
        RECT 12.535 181.340 14.495 181.570 ;
        RECT 15.215 180.880 16.545 190.670 ;
        RECT 45.135 190.570 49.450 190.670 ;
        RECT 56.110 190.570 56.570 207.460 ;
        RECT 17.265 189.980 19.225 190.210 ;
        RECT 19.555 189.980 21.515 190.210 ;
        RECT 21.845 189.980 23.805 190.210 ;
        RECT 24.135 189.980 26.095 190.210 ;
        RECT 26.425 189.980 28.385 190.210 ;
        RECT 28.715 189.980 30.675 190.210 ;
        RECT 31.005 189.980 32.965 190.210 ;
        RECT 33.295 189.980 35.255 190.210 ;
        RECT 35.585 189.980 37.545 190.210 ;
        RECT 37.875 189.980 39.835 190.210 ;
        RECT 40.165 189.980 42.125 190.210 ;
        RECT 42.455 189.980 44.415 190.210 ;
        RECT 16.985 189.645 17.215 189.775 ;
        RECT 16.950 188.245 17.250 189.645 ;
        RECT 16.985 181.775 17.215 188.245 ;
        RECT 19.275 186.555 19.505 189.775 ;
        RECT 21.565 189.645 21.795 189.775 ;
        RECT 21.530 188.245 21.830 189.645 ;
        RECT 19.240 184.995 19.540 186.555 ;
        RECT 19.275 181.775 19.505 184.995 ;
        RECT 21.565 181.775 21.795 188.245 ;
        RECT 23.855 186.555 24.085 189.775 ;
        RECT 26.145 189.645 26.375 189.775 ;
        RECT 26.110 188.245 26.410 189.645 ;
        RECT 23.820 184.995 24.120 186.555 ;
        RECT 23.855 181.775 24.085 184.995 ;
        RECT 26.145 181.775 26.375 188.245 ;
        RECT 28.435 186.555 28.665 189.775 ;
        RECT 30.725 189.645 30.955 189.775 ;
        RECT 30.690 188.245 30.990 189.645 ;
        RECT 28.400 184.995 28.700 186.555 ;
        RECT 28.435 181.775 28.665 184.995 ;
        RECT 30.725 181.775 30.955 188.245 ;
        RECT 33.015 186.555 33.245 189.775 ;
        RECT 35.305 189.645 35.535 189.775 ;
        RECT 35.270 188.245 35.570 189.645 ;
        RECT 32.980 184.995 33.280 186.555 ;
        RECT 33.015 181.775 33.245 184.995 ;
        RECT 35.305 181.775 35.535 188.245 ;
        RECT 37.595 186.555 37.825 189.775 ;
        RECT 39.885 189.645 40.115 189.775 ;
        RECT 39.850 188.245 40.150 189.645 ;
        RECT 37.560 184.995 37.860 186.555 ;
        RECT 37.595 181.775 37.825 184.995 ;
        RECT 39.885 181.775 40.115 188.245 ;
        RECT 42.175 186.555 42.405 189.775 ;
        RECT 44.465 189.645 44.695 189.775 ;
        RECT 44.430 188.245 44.730 189.645 ;
        RECT 42.140 184.995 42.440 186.555 ;
        RECT 42.175 181.775 42.405 184.995 ;
        RECT 44.465 181.775 44.695 188.245 ;
        RECT 45.135 187.880 50.745 190.570 ;
        RECT 51.315 188.465 53.075 190.570 ;
        RECT 53.655 188.465 54.245 190.570 ;
        RECT 54.825 188.465 56.570 190.570 ;
        RECT 54.835 187.880 56.570 188.465 ;
        RECT 45.135 187.650 56.570 187.880 ;
        RECT 17.465 181.570 19.025 181.605 ;
        RECT 19.755 181.570 21.315 181.605 ;
        RECT 22.045 181.570 23.605 181.605 ;
        RECT 24.335 181.570 25.895 181.605 ;
        RECT 26.625 181.570 28.185 181.605 ;
        RECT 28.915 181.570 30.475 181.605 ;
        RECT 31.205 181.570 32.765 181.605 ;
        RECT 33.495 181.570 35.055 181.605 ;
        RECT 35.785 181.570 37.345 181.605 ;
        RECT 38.075 181.570 39.635 181.605 ;
        RECT 40.365 181.570 41.925 181.605 ;
        RECT 42.655 181.570 44.215 181.605 ;
        RECT 17.265 181.340 44.415 181.570 ;
        RECT 17.465 181.305 19.025 181.340 ;
        RECT 19.755 181.305 21.315 181.340 ;
        RECT 22.045 181.305 23.605 181.340 ;
        RECT 24.335 181.305 25.895 181.340 ;
        RECT 26.625 181.305 28.185 181.340 ;
        RECT 28.915 181.305 30.475 181.340 ;
        RECT 31.205 181.305 32.765 181.340 ;
        RECT 33.495 181.305 35.055 181.340 ;
        RECT 35.785 181.305 37.345 181.340 ;
        RECT 38.075 181.305 39.635 181.340 ;
        RECT 40.365 181.305 41.925 181.340 ;
        RECT 42.655 181.305 44.215 181.340 ;
        RECT 45.135 180.880 46.085 187.650 ;
        RECT 4.100 180.050 46.085 180.880 ;
        RECT 4.100 127.485 4.900 180.050 ;
        RECT 5.910 178.420 53.180 179.250 ;
        RECT 5.910 168.720 9.530 178.420 ;
        RECT 17.400 177.960 18.800 178.130 ;
        RECT 19.690 177.960 21.090 178.130 ;
        RECT 26.560 177.960 27.960 178.130 ;
        RECT 28.850 177.960 30.250 178.130 ;
        RECT 35.720 177.960 37.120 178.130 ;
        RECT 38.010 177.960 39.410 178.130 ;
        RECT 44.880 177.960 46.280 178.130 ;
        RECT 47.170 177.960 48.570 178.130 ;
        RECT 49.460 177.960 50.860 178.130 ;
        RECT 10.250 177.730 12.210 177.960 ;
        RECT 12.540 177.730 14.500 177.960 ;
        RECT 14.830 177.730 16.790 177.960 ;
        RECT 17.120 177.730 19.080 177.960 ;
        RECT 19.410 177.730 21.370 177.960 ;
        RECT 21.700 177.730 23.660 177.960 ;
        RECT 23.990 177.730 25.950 177.960 ;
        RECT 26.280 177.730 28.240 177.960 ;
        RECT 28.570 177.730 30.530 177.960 ;
        RECT 30.860 177.730 32.820 177.960 ;
        RECT 33.150 177.730 35.110 177.960 ;
        RECT 35.440 177.730 37.400 177.960 ;
        RECT 37.730 177.730 39.690 177.960 ;
        RECT 40.020 177.730 41.980 177.960 ;
        RECT 42.310 177.730 44.270 177.960 ;
        RECT 44.600 177.730 46.560 177.960 ;
        RECT 46.890 177.730 48.850 177.960 ;
        RECT 49.180 177.730 51.140 177.960 ;
        RECT 9.970 174.270 10.200 177.570 ;
        RECT 12.260 174.270 12.490 177.570 ;
        RECT 14.550 176.670 14.780 177.570 ;
        RECT 14.465 175.270 14.865 176.670 ;
        RECT 9.885 172.870 10.285 174.270 ;
        RECT 12.175 172.870 12.575 174.270 ;
        RECT 9.970 169.570 10.200 172.870 ;
        RECT 12.260 169.570 12.490 172.870 ;
        RECT 14.550 169.570 14.780 175.270 ;
        RECT 16.840 174.270 17.070 177.570 ;
        RECT 16.755 172.870 17.155 174.270 ;
        RECT 16.840 169.570 17.070 172.870 ;
        RECT 19.130 171.870 19.360 177.570 ;
        RECT 21.420 174.270 21.650 177.570 ;
        RECT 23.710 176.670 23.940 177.570 ;
        RECT 23.625 175.270 24.025 176.670 ;
        RECT 21.335 172.870 21.735 174.270 ;
        RECT 19.045 170.470 19.445 171.870 ;
        RECT 19.130 169.570 19.360 170.470 ;
        RECT 21.420 169.570 21.650 172.870 ;
        RECT 23.710 169.570 23.940 175.270 ;
        RECT 26.000 174.270 26.230 177.570 ;
        RECT 25.915 172.870 26.315 174.270 ;
        RECT 26.000 169.570 26.230 172.870 ;
        RECT 28.290 171.870 28.520 177.570 ;
        RECT 30.580 174.270 30.810 177.570 ;
        RECT 32.870 176.670 33.100 177.570 ;
        RECT 32.785 175.270 33.185 176.670 ;
        RECT 30.495 172.870 30.895 174.270 ;
        RECT 28.205 170.470 28.605 171.870 ;
        RECT 28.290 169.570 28.520 170.470 ;
        RECT 30.580 169.570 30.810 172.870 ;
        RECT 32.870 169.570 33.100 175.270 ;
        RECT 35.160 174.270 35.390 177.570 ;
        RECT 35.075 172.870 35.475 174.270 ;
        RECT 35.160 169.570 35.390 172.870 ;
        RECT 37.450 171.870 37.680 177.570 ;
        RECT 39.740 174.270 39.970 177.570 ;
        RECT 42.030 176.670 42.260 177.570 ;
        RECT 41.945 175.270 42.345 176.670 ;
        RECT 39.655 172.870 40.055 174.270 ;
        RECT 37.365 170.470 37.765 171.870 ;
        RECT 37.450 169.570 37.680 170.470 ;
        RECT 39.740 169.570 39.970 172.870 ;
        RECT 42.030 169.570 42.260 175.270 ;
        RECT 44.320 174.270 44.550 177.570 ;
        RECT 44.235 172.870 44.635 174.270 ;
        RECT 44.320 169.570 44.550 172.870 ;
        RECT 46.610 171.870 46.840 177.570 ;
        RECT 48.900 174.270 49.130 177.570 ;
        RECT 51.190 174.270 51.420 177.570 ;
        RECT 48.815 172.870 49.215 174.270 ;
        RECT 51.105 172.870 51.505 174.270 ;
        RECT 46.525 170.470 46.925 171.870 ;
        RECT 46.610 169.570 46.840 170.470 ;
        RECT 48.900 169.570 49.130 172.870 ;
        RECT 51.190 169.570 51.420 172.870 ;
        RECT 10.250 169.180 12.210 169.410 ;
        RECT 12.540 169.180 14.500 169.410 ;
        RECT 14.830 169.180 16.790 169.410 ;
        RECT 17.120 169.180 19.080 169.410 ;
        RECT 19.410 169.180 21.370 169.410 ;
        RECT 21.700 169.180 23.660 169.410 ;
        RECT 23.990 169.180 25.950 169.410 ;
        RECT 26.280 169.180 28.240 169.410 ;
        RECT 28.570 169.180 30.530 169.410 ;
        RECT 30.860 169.180 32.820 169.410 ;
        RECT 33.150 169.180 35.110 169.410 ;
        RECT 35.440 169.180 37.400 169.410 ;
        RECT 37.730 169.180 39.690 169.410 ;
        RECT 40.020 169.180 41.980 169.410 ;
        RECT 42.310 169.180 44.270 169.410 ;
        RECT 44.600 169.180 46.560 169.410 ;
        RECT 46.890 169.180 48.850 169.410 ;
        RECT 49.180 169.180 51.140 169.410 ;
        RECT 10.530 169.010 11.930 169.180 ;
        RECT 12.820 169.010 14.220 169.180 ;
        RECT 15.110 169.010 16.510 169.180 ;
        RECT 21.980 169.010 23.380 169.180 ;
        RECT 24.270 169.010 25.670 169.180 ;
        RECT 31.140 169.010 32.540 169.180 ;
        RECT 33.430 169.010 34.830 169.180 ;
        RECT 40.300 169.010 41.700 169.180 ;
        RECT 42.590 169.010 43.990 169.180 ;
        RECT 51.860 168.720 53.180 178.420 ;
        RECT 5.910 167.830 53.180 168.720 ;
        RECT 5.910 148.290 9.530 167.830 ;
        RECT 10.310 167.140 12.270 167.370 ;
        RECT 12.600 167.140 14.560 167.370 ;
        RECT 16.350 167.140 18.310 167.370 ;
        RECT 18.640 167.140 20.600 167.370 ;
        RECT 22.390 167.140 24.350 167.370 ;
        RECT 24.680 167.140 26.640 167.370 ;
        RECT 28.430 167.140 30.390 167.370 ;
        RECT 30.720 167.140 32.680 167.370 ;
        RECT 34.470 167.140 36.430 167.370 ;
        RECT 36.760 167.140 38.720 167.370 ;
        RECT 40.510 167.140 42.470 167.370 ;
        RECT 42.800 167.140 44.760 167.370 ;
        RECT 46.550 167.140 48.510 167.370 ;
        RECT 48.840 167.140 50.800 167.370 ;
        RECT 10.030 161.265 10.260 166.980 ;
        RECT 12.320 161.265 12.550 166.980 ;
        RECT 14.610 161.265 14.840 166.980 ;
        RECT 16.070 161.265 16.300 166.980 ;
        RECT 18.360 166.565 18.590 166.980 ;
        RECT 18.325 165.865 18.625 166.565 ;
        RECT 9.995 159.865 10.295 161.265 ;
        RECT 12.285 159.865 12.585 161.265 ;
        RECT 14.575 159.865 14.875 161.265 ;
        RECT 16.035 159.865 16.335 161.265 ;
        RECT 10.030 158.820 10.260 159.865 ;
        RECT 12.320 158.820 12.550 159.865 ;
        RECT 14.610 158.820 14.840 159.865 ;
        RECT 16.070 158.980 16.300 159.865 ;
        RECT 18.360 158.980 18.590 165.865 ;
        RECT 20.650 161.265 20.880 166.980 ;
        RECT 22.110 161.265 22.340 166.980 ;
        RECT 24.400 166.565 24.630 166.980 ;
        RECT 24.365 165.865 24.665 166.565 ;
        RECT 20.615 159.865 20.915 161.265 ;
        RECT 22.075 159.865 22.375 161.265 ;
        RECT 20.650 158.980 20.880 159.865 ;
        RECT 22.110 158.980 22.340 159.865 ;
        RECT 24.400 158.980 24.630 165.865 ;
        RECT 26.690 161.265 26.920 166.980 ;
        RECT 28.150 161.265 28.380 166.980 ;
        RECT 30.440 162.965 30.670 166.980 ;
        RECT 30.405 162.265 30.705 162.965 ;
        RECT 26.655 159.865 26.955 161.265 ;
        RECT 28.115 159.865 28.415 161.265 ;
        RECT 26.690 158.980 26.920 159.865 ;
        RECT 28.150 158.980 28.380 159.865 ;
        RECT 30.440 158.980 30.670 162.265 ;
        RECT 32.730 161.265 32.960 166.980 ;
        RECT 34.190 161.265 34.420 166.980 ;
        RECT 36.480 166.565 36.710 166.980 ;
        RECT 36.445 165.865 36.745 166.565 ;
        RECT 32.695 159.865 32.995 161.265 ;
        RECT 34.155 159.865 34.455 161.265 ;
        RECT 32.730 158.980 32.960 159.865 ;
        RECT 34.190 158.980 34.420 159.865 ;
        RECT 36.480 158.980 36.710 165.865 ;
        RECT 38.770 161.265 39.000 166.980 ;
        RECT 40.230 161.265 40.460 166.980 ;
        RECT 42.520 166.565 42.750 166.980 ;
        RECT 42.485 165.865 42.785 166.565 ;
        RECT 38.735 159.865 39.035 161.265 ;
        RECT 40.195 159.865 40.495 161.265 ;
        RECT 38.770 158.980 39.000 159.865 ;
        RECT 40.230 158.980 40.460 159.865 ;
        RECT 42.520 158.980 42.750 165.865 ;
        RECT 44.810 161.265 45.040 166.980 ;
        RECT 46.270 161.265 46.500 166.980 ;
        RECT 48.560 161.265 48.790 166.980 ;
        RECT 50.850 161.265 51.080 166.980 ;
        RECT 44.775 159.865 45.075 161.265 ;
        RECT 46.235 159.865 46.535 161.265 ;
        RECT 48.525 159.865 48.825 161.265 ;
        RECT 50.815 159.865 51.115 161.265 ;
        RECT 44.810 158.980 45.040 159.865 ;
        RECT 46.270 158.820 46.500 159.865 ;
        RECT 48.560 158.820 48.790 159.865 ;
        RECT 50.850 158.820 51.080 159.865 ;
        RECT 10.030 158.590 14.840 158.820 ;
        RECT 10.030 157.210 14.840 157.440 ;
        RECT 16.350 157.210 44.760 158.820 ;
        RECT 46.270 158.590 51.080 158.820 ;
        RECT 46.270 157.210 51.080 157.440 ;
        RECT 10.030 156.165 10.260 157.210 ;
        RECT 12.320 156.165 12.550 157.210 ;
        RECT 14.610 156.165 14.840 157.210 ;
        RECT 16.070 156.165 16.300 157.050 ;
        RECT 9.995 154.765 10.295 156.165 ;
        RECT 12.285 154.765 12.585 156.165 ;
        RECT 14.575 154.765 14.875 156.165 ;
        RECT 16.035 154.765 16.335 156.165 ;
        RECT 10.030 149.050 10.260 154.765 ;
        RECT 12.320 149.050 12.550 154.765 ;
        RECT 14.610 149.050 14.840 154.765 ;
        RECT 16.070 149.050 16.300 154.765 ;
        RECT 18.360 150.165 18.590 157.050 ;
        RECT 20.650 156.165 20.880 157.050 ;
        RECT 22.110 156.165 22.340 157.050 ;
        RECT 20.615 154.765 20.915 156.165 ;
        RECT 22.075 154.765 22.375 156.165 ;
        RECT 18.325 149.465 18.625 150.165 ;
        RECT 18.360 149.050 18.590 149.465 ;
        RECT 20.650 149.050 20.880 154.765 ;
        RECT 22.110 149.050 22.340 154.765 ;
        RECT 24.400 151.965 24.630 157.050 ;
        RECT 26.690 156.165 26.920 157.050 ;
        RECT 28.150 156.165 28.380 157.050 ;
        RECT 26.655 154.765 26.955 156.165 ;
        RECT 28.115 154.765 28.415 156.165 ;
        RECT 24.365 151.265 24.665 151.965 ;
        RECT 24.400 149.050 24.630 151.265 ;
        RECT 26.690 149.050 26.920 154.765 ;
        RECT 28.150 149.050 28.380 154.765 ;
        RECT 30.440 149.050 30.670 157.210 ;
        RECT 32.730 156.165 32.960 157.050 ;
        RECT 32.695 154.765 32.995 156.165 ;
        RECT 32.730 149.050 32.960 154.765 ;
        RECT 34.190 149.050 34.420 157.210 ;
        RECT 36.480 149.050 36.710 157.210 ;
        RECT 38.770 149.050 39.000 157.210 ;
        RECT 40.230 156.165 40.460 157.050 ;
        RECT 40.195 154.765 40.495 156.165 ;
        RECT 40.230 149.050 40.460 154.765 ;
        RECT 42.520 150.165 42.750 157.050 ;
        RECT 44.810 156.165 45.040 157.050 ;
        RECT 46.270 156.165 46.500 157.210 ;
        RECT 48.560 156.165 48.790 157.210 ;
        RECT 50.850 156.165 51.080 157.210 ;
        RECT 44.775 154.765 45.075 156.165 ;
        RECT 46.235 154.765 46.535 156.165 ;
        RECT 48.525 154.765 48.825 156.165 ;
        RECT 50.815 154.765 51.115 156.165 ;
        RECT 42.485 149.465 42.785 150.165 ;
        RECT 42.520 149.050 42.750 149.465 ;
        RECT 44.810 149.050 45.040 154.765 ;
        RECT 46.270 149.050 46.500 154.765 ;
        RECT 48.560 149.050 48.790 154.765 ;
        RECT 50.850 149.050 51.080 154.765 ;
        RECT 10.310 148.660 12.270 148.890 ;
        RECT 12.600 148.660 14.560 148.890 ;
        RECT 16.350 148.660 18.310 148.890 ;
        RECT 18.640 148.660 20.600 148.890 ;
        RECT 22.390 148.660 24.350 148.890 ;
        RECT 24.680 148.660 26.640 148.890 ;
        RECT 28.430 148.660 30.390 148.890 ;
        RECT 30.720 148.660 32.680 148.890 ;
        RECT 34.470 148.660 36.430 148.890 ;
        RECT 36.760 148.660 38.720 148.890 ;
        RECT 40.510 148.660 42.470 148.890 ;
        RECT 42.800 148.660 44.760 148.890 ;
        RECT 46.550 148.660 48.510 148.890 ;
        RECT 48.840 148.660 50.800 148.890 ;
        RECT 51.580 148.290 53.180 167.830 ;
        RECT 5.910 143.745 53.180 148.290 ;
        RECT 62.865 171.445 63.455 212.490 ;
        RECT 63.895 211.600 64.595 212.600 ;
        RECT 77.595 212.570 78.595 212.805 ;
        RECT 77.595 211.395 78.595 211.630 ;
        RECT 80.185 211.600 81.755 212.600 ;
        RECT 83.345 212.570 84.345 212.805 ;
        RECT 83.345 211.395 84.345 211.630 ;
        RECT 97.345 211.600 98.045 212.600 ;
        RECT 64.175 211.165 80.135 211.395 ;
        RECT 81.805 211.165 97.765 211.395 ;
        RECT 77.595 210.930 78.595 211.165 ;
        RECT 83.345 210.930 84.345 211.165 ;
        RECT 77.595 210.015 78.595 210.250 ;
        RECT 83.345 210.015 84.345 210.250 ;
        RECT 64.175 209.785 80.135 210.015 ;
        RECT 81.805 209.785 97.765 210.015 ;
        RECT 63.895 208.580 64.595 209.580 ;
        RECT 77.595 209.550 78.595 209.785 ;
        RECT 77.595 208.375 78.595 208.610 ;
        RECT 80.185 208.580 81.755 209.580 ;
        RECT 83.345 209.550 84.345 209.785 ;
        RECT 83.345 208.375 84.345 208.610 ;
        RECT 97.345 208.580 98.045 209.580 ;
        RECT 64.175 208.145 80.135 208.375 ;
        RECT 81.805 208.145 97.765 208.375 ;
        RECT 77.595 207.910 78.595 208.145 ;
        RECT 83.345 207.910 84.345 208.145 ;
        RECT 77.595 206.995 78.595 207.230 ;
        RECT 83.345 206.995 84.345 207.230 ;
        RECT 64.175 206.765 80.135 206.995 ;
        RECT 81.805 206.765 97.765 206.995 ;
        RECT 63.895 205.560 64.595 206.560 ;
        RECT 77.595 206.530 78.595 206.765 ;
        RECT 77.595 205.355 78.595 205.590 ;
        RECT 80.185 205.560 81.755 206.560 ;
        RECT 83.345 206.530 84.345 206.765 ;
        RECT 83.345 205.355 84.345 205.590 ;
        RECT 97.345 205.560 98.045 206.560 ;
        RECT 64.175 205.125 80.135 205.355 ;
        RECT 81.805 205.125 97.765 205.355 ;
        RECT 77.595 204.890 78.595 205.125 ;
        RECT 83.345 204.890 84.345 205.125 ;
        RECT 77.595 203.975 78.595 204.210 ;
        RECT 83.345 203.975 84.345 204.210 ;
        RECT 64.175 203.745 80.135 203.975 ;
        RECT 81.805 203.745 97.765 203.975 ;
        RECT 63.895 202.540 75.695 203.540 ;
        RECT 77.595 203.510 78.595 203.745 ;
        RECT 77.595 202.335 78.595 202.570 ;
        RECT 80.185 202.540 81.755 203.540 ;
        RECT 83.345 203.510 84.345 203.745 ;
        RECT 83.345 202.335 84.345 202.570 ;
        RECT 86.245 202.540 98.045 203.540 ;
        RECT 64.175 202.105 80.135 202.335 ;
        RECT 81.805 202.105 97.765 202.335 ;
        RECT 77.595 201.870 78.595 202.105 ;
        RECT 83.345 201.870 84.345 202.105 ;
        RECT 77.595 200.955 78.595 201.190 ;
        RECT 83.345 200.955 84.345 201.190 ;
        RECT 64.175 200.725 80.135 200.955 ;
        RECT 81.805 200.725 97.765 200.955 ;
        RECT 63.895 199.520 70.195 200.520 ;
        RECT 77.595 200.490 78.595 200.725 ;
        RECT 77.595 199.315 78.595 199.550 ;
        RECT 80.185 199.520 81.755 200.520 ;
        RECT 83.345 200.490 84.345 200.725 ;
        RECT 83.345 199.315 84.345 199.550 ;
        RECT 91.745 199.520 98.045 200.520 ;
        RECT 64.175 199.085 80.135 199.315 ;
        RECT 81.805 199.085 97.765 199.315 ;
        RECT 77.595 198.850 78.595 199.085 ;
        RECT 83.345 198.850 84.345 199.085 ;
        RECT 77.595 197.935 78.595 198.170 ;
        RECT 83.345 197.935 84.345 198.170 ;
        RECT 64.175 197.705 80.135 197.935 ;
        RECT 81.805 197.705 97.765 197.935 ;
        RECT 63.895 196.500 67.445 197.500 ;
        RECT 77.595 197.470 78.595 197.705 ;
        RECT 77.595 196.295 78.595 196.530 ;
        RECT 80.185 196.500 81.755 197.500 ;
        RECT 83.345 197.470 84.345 197.705 ;
        RECT 83.345 196.295 84.345 196.530 ;
        RECT 94.495 196.500 98.045 197.500 ;
        RECT 64.175 196.065 80.135 196.295 ;
        RECT 81.805 196.065 97.765 196.295 ;
        RECT 77.595 195.830 78.595 196.065 ;
        RECT 83.345 195.830 84.345 196.065 ;
        RECT 77.595 194.915 78.595 195.150 ;
        RECT 83.345 194.915 84.345 195.150 ;
        RECT 64.175 194.685 80.135 194.915 ;
        RECT 81.805 194.685 97.765 194.915 ;
        RECT 63.895 193.480 72.945 194.480 ;
        RECT 77.595 194.450 78.595 194.685 ;
        RECT 77.595 193.275 78.595 193.510 ;
        RECT 80.185 193.480 81.755 194.480 ;
        RECT 83.345 194.450 84.345 194.685 ;
        RECT 83.345 193.275 84.345 193.510 ;
        RECT 88.995 193.480 98.045 194.480 ;
        RECT 64.175 193.045 80.135 193.275 ;
        RECT 81.805 193.045 97.765 193.275 ;
        RECT 77.595 192.810 78.595 193.045 ;
        RECT 83.345 192.810 84.345 193.045 ;
        RECT 77.595 191.895 78.595 192.130 ;
        RECT 83.345 191.895 84.345 192.130 ;
        RECT 64.175 191.665 80.135 191.895 ;
        RECT 81.805 191.665 97.765 191.895 ;
        RECT 63.895 190.460 67.445 191.460 ;
        RECT 77.595 191.430 78.595 191.665 ;
        RECT 77.595 190.255 78.595 190.490 ;
        RECT 80.185 190.460 81.755 191.460 ;
        RECT 83.345 191.430 84.345 191.665 ;
        RECT 83.345 190.255 84.345 190.490 ;
        RECT 94.495 190.460 98.045 191.460 ;
        RECT 64.175 190.025 80.135 190.255 ;
        RECT 81.805 190.025 97.765 190.255 ;
        RECT 77.595 189.790 78.595 190.025 ;
        RECT 83.345 189.790 84.345 190.025 ;
        RECT 77.595 188.875 78.595 189.110 ;
        RECT 83.345 188.875 84.345 189.110 ;
        RECT 64.175 188.645 80.135 188.875 ;
        RECT 81.805 188.645 97.765 188.875 ;
        RECT 63.895 187.440 70.195 188.440 ;
        RECT 77.595 188.410 78.595 188.645 ;
        RECT 77.595 187.235 78.595 187.470 ;
        RECT 80.185 187.440 81.755 188.440 ;
        RECT 83.345 188.410 84.345 188.645 ;
        RECT 83.345 187.235 84.345 187.470 ;
        RECT 91.745 187.440 98.045 188.440 ;
        RECT 64.175 187.005 80.135 187.235 ;
        RECT 81.805 187.005 97.765 187.235 ;
        RECT 77.595 186.770 78.595 187.005 ;
        RECT 83.345 186.770 84.345 187.005 ;
        RECT 77.595 185.855 78.595 186.090 ;
        RECT 83.345 185.855 84.345 186.090 ;
        RECT 64.175 185.625 80.135 185.855 ;
        RECT 81.805 185.625 97.765 185.855 ;
        RECT 63.895 184.420 75.695 185.420 ;
        RECT 77.595 185.390 78.595 185.625 ;
        RECT 77.595 184.215 78.595 184.450 ;
        RECT 80.185 184.420 81.755 185.420 ;
        RECT 83.345 185.390 84.345 185.625 ;
        RECT 83.345 184.215 84.345 184.450 ;
        RECT 86.245 184.420 98.045 185.420 ;
        RECT 64.175 183.985 80.135 184.215 ;
        RECT 81.805 183.985 97.765 184.215 ;
        RECT 77.595 183.750 78.595 183.985 ;
        RECT 83.345 183.750 84.345 183.985 ;
        RECT 77.595 182.835 78.595 183.070 ;
        RECT 83.345 182.835 84.345 183.070 ;
        RECT 64.175 182.605 80.135 182.835 ;
        RECT 81.805 182.605 97.765 182.835 ;
        RECT 98.485 182.710 102.825 216.515 ;
        RECT 108.520 216.690 108.920 217.515 ;
        RECT 109.325 217.500 109.555 217.755 ;
        RECT 110.615 217.500 110.845 217.755 ;
        RECT 111.905 217.500 112.135 217.755 ;
        RECT 109.605 216.945 110.565 217.295 ;
        RECT 110.895 217.065 111.855 217.295 ;
        RECT 112.545 216.690 112.950 220.315 ;
        RECT 113.635 219.705 114.595 219.935 ;
        RECT 114.925 219.705 115.885 220.055 ;
        RECT 113.355 219.255 113.585 219.500 ;
        RECT 114.645 219.255 114.875 219.500 ;
        RECT 115.935 219.255 116.165 219.500 ;
        RECT 113.320 217.755 113.620 219.255 ;
        RECT 114.610 217.755 114.910 219.255 ;
        RECT 115.900 217.755 116.200 219.255 ;
        RECT 113.355 217.500 113.585 217.755 ;
        RECT 114.645 217.500 114.875 217.755 ;
        RECT 115.935 217.500 116.165 217.755 ;
        RECT 113.635 216.945 114.595 217.295 ;
        RECT 114.925 217.065 115.885 217.295 ;
        RECT 116.575 216.690 116.980 220.315 ;
        RECT 117.665 219.705 118.625 219.935 ;
        RECT 118.955 219.705 119.915 220.055 ;
        RECT 117.385 219.255 117.615 219.500 ;
        RECT 118.675 219.255 118.905 219.500 ;
        RECT 119.965 219.255 120.195 219.500 ;
        RECT 117.350 217.755 117.650 219.255 ;
        RECT 118.640 217.755 118.940 219.255 ;
        RECT 119.930 217.755 120.230 219.255 ;
        RECT 117.385 217.500 117.615 217.755 ;
        RECT 118.675 217.500 118.905 217.755 ;
        RECT 119.965 217.500 120.195 217.755 ;
        RECT 117.665 216.945 118.625 217.295 ;
        RECT 118.955 217.065 119.915 217.295 ;
        RECT 120.605 216.690 121.010 220.315 ;
        RECT 121.695 219.705 122.655 219.935 ;
        RECT 122.985 219.705 123.945 220.055 ;
        RECT 121.415 219.255 121.645 219.500 ;
        RECT 122.705 219.255 122.935 219.500 ;
        RECT 123.995 219.255 124.225 219.500 ;
        RECT 121.380 217.755 121.680 219.255 ;
        RECT 122.670 217.755 122.970 219.255 ;
        RECT 123.960 217.755 124.260 219.255 ;
        RECT 121.415 217.500 121.645 217.755 ;
        RECT 122.705 217.500 122.935 217.755 ;
        RECT 123.995 217.500 124.225 217.755 ;
        RECT 121.695 216.945 122.655 217.295 ;
        RECT 122.985 217.065 123.945 217.295 ;
        RECT 124.635 216.690 125.040 220.315 ;
        RECT 125.725 219.705 126.685 219.935 ;
        RECT 127.015 219.705 127.975 220.055 ;
        RECT 125.445 219.255 125.675 219.500 ;
        RECT 126.735 219.255 126.965 219.500 ;
        RECT 128.025 219.255 128.255 219.500 ;
        RECT 125.410 217.755 125.710 219.255 ;
        RECT 126.700 217.755 127.000 219.255 ;
        RECT 127.990 217.755 128.290 219.255 ;
        RECT 125.445 217.500 125.675 217.755 ;
        RECT 126.735 217.500 126.965 217.755 ;
        RECT 128.025 217.500 128.255 217.755 ;
        RECT 125.725 216.945 126.685 217.295 ;
        RECT 127.015 217.065 127.975 217.295 ;
        RECT 128.665 216.690 129.070 220.315 ;
        RECT 129.755 219.705 130.715 219.935 ;
        RECT 131.045 219.705 132.005 220.055 ;
        RECT 129.475 219.255 129.705 219.500 ;
        RECT 130.765 219.255 130.995 219.500 ;
        RECT 132.055 219.255 132.285 219.500 ;
        RECT 129.440 217.755 129.740 219.255 ;
        RECT 130.730 217.755 131.030 219.255 ;
        RECT 132.020 217.755 132.320 219.255 ;
        RECT 129.475 217.500 129.705 217.755 ;
        RECT 130.765 217.500 130.995 217.755 ;
        RECT 132.055 217.500 132.285 217.755 ;
        RECT 129.755 216.945 130.715 217.295 ;
        RECT 131.045 217.065 132.005 217.295 ;
        RECT 132.695 216.690 133.100 220.315 ;
        RECT 133.785 219.705 134.745 219.935 ;
        RECT 135.075 219.705 136.035 220.055 ;
        RECT 133.505 219.255 133.735 219.500 ;
        RECT 134.795 219.255 135.025 219.500 ;
        RECT 136.085 219.255 136.315 219.500 ;
        RECT 133.470 217.755 133.770 219.255 ;
        RECT 134.760 217.755 135.060 219.255 ;
        RECT 136.050 217.755 136.350 219.255 ;
        RECT 133.505 217.500 133.735 217.755 ;
        RECT 134.795 217.500 135.025 217.755 ;
        RECT 136.085 217.500 136.315 217.755 ;
        RECT 133.785 216.945 134.745 217.295 ;
        RECT 135.075 217.065 136.035 217.295 ;
        RECT 136.725 216.690 137.130 220.315 ;
        RECT 137.815 219.705 138.775 219.935 ;
        RECT 139.105 219.705 140.065 220.055 ;
        RECT 137.535 219.255 137.765 219.500 ;
        RECT 138.825 219.255 139.055 219.500 ;
        RECT 140.115 219.255 140.345 219.500 ;
        RECT 137.500 217.755 137.800 219.255 ;
        RECT 138.790 217.755 139.090 219.255 ;
        RECT 140.080 217.755 140.380 219.255 ;
        RECT 137.535 217.500 137.765 217.755 ;
        RECT 138.825 217.500 139.055 217.755 ;
        RECT 140.115 217.500 140.345 217.755 ;
        RECT 137.815 216.945 138.775 217.295 ;
        RECT 139.105 217.065 140.065 217.295 ;
        RECT 140.755 216.690 141.160 220.315 ;
        RECT 141.845 219.705 142.805 219.935 ;
        RECT 143.135 219.705 144.095 220.055 ;
        RECT 141.565 219.255 141.795 219.500 ;
        RECT 142.855 219.255 143.085 219.500 ;
        RECT 144.145 219.255 144.375 219.500 ;
        RECT 141.530 217.755 141.830 219.255 ;
        RECT 142.820 217.755 143.120 219.255 ;
        RECT 144.110 217.755 144.410 219.255 ;
        RECT 141.565 217.500 141.795 217.755 ;
        RECT 142.855 217.500 143.085 217.755 ;
        RECT 144.145 217.500 144.375 217.755 ;
        RECT 141.845 216.945 142.805 217.295 ;
        RECT 143.135 217.065 144.095 217.295 ;
        RECT 144.785 216.690 145.190 220.315 ;
        RECT 145.875 219.705 146.835 219.935 ;
        RECT 147.165 219.705 148.125 220.055 ;
        RECT 145.595 219.255 145.825 219.500 ;
        RECT 146.885 219.255 147.115 219.500 ;
        RECT 148.175 219.255 148.405 219.500 ;
        RECT 145.560 217.755 145.860 219.255 ;
        RECT 146.850 217.755 147.150 219.255 ;
        RECT 148.140 217.755 148.440 219.255 ;
        RECT 145.595 217.500 145.825 217.755 ;
        RECT 146.885 217.500 147.115 217.755 ;
        RECT 148.175 217.500 148.405 217.755 ;
        RECT 145.875 216.945 146.835 217.295 ;
        RECT 147.165 217.065 148.125 217.295 ;
        RECT 148.815 216.690 149.220 220.315 ;
        RECT 149.905 219.705 150.865 219.935 ;
        RECT 151.195 219.705 152.155 220.055 ;
        RECT 149.625 219.255 149.855 219.500 ;
        RECT 150.915 219.255 151.145 219.500 ;
        RECT 152.205 219.255 152.435 219.500 ;
        RECT 149.590 217.755 149.890 219.255 ;
        RECT 150.880 217.755 151.180 219.255 ;
        RECT 152.170 217.755 152.470 219.255 ;
        RECT 149.625 217.500 149.855 217.755 ;
        RECT 150.915 217.500 151.145 217.755 ;
        RECT 152.205 217.500 152.435 217.755 ;
        RECT 149.905 216.945 150.865 217.295 ;
        RECT 151.195 217.065 152.155 217.295 ;
        RECT 152.845 216.690 153.245 220.315 ;
        RECT 108.520 216.290 153.245 216.690 ;
        RECT 106.415 213.340 153.245 213.740 ;
        RECT 106.415 210.540 108.915 213.340 ;
        RECT 109.605 212.735 110.565 212.965 ;
        RECT 110.895 212.735 111.855 212.965 ;
        RECT 108.515 203.720 108.915 210.540 ;
        RECT 109.325 205.495 109.555 212.530 ;
        RECT 110.615 211.190 110.845 212.530 ;
        RECT 110.580 209.690 110.880 211.190 ;
        RECT 109.290 204.795 109.590 205.495 ;
        RECT 109.325 204.530 109.555 204.795 ;
        RECT 110.615 204.530 110.845 209.690 ;
        RECT 111.905 206.705 112.135 212.530 ;
        RECT 111.870 206.005 112.170 206.705 ;
        RECT 111.905 204.530 112.135 206.005 ;
        RECT 109.605 203.995 110.565 204.325 ;
        RECT 110.895 203.995 111.855 204.325 ;
        RECT 112.545 203.720 112.945 213.340 ;
        RECT 113.635 212.735 114.595 212.965 ;
        RECT 114.925 212.735 115.885 212.965 ;
        RECT 113.355 205.495 113.585 212.530 ;
        RECT 114.645 211.190 114.875 212.530 ;
        RECT 114.610 209.690 114.910 211.190 ;
        RECT 113.320 204.795 113.620 205.495 ;
        RECT 113.355 204.530 113.585 204.795 ;
        RECT 114.645 204.530 114.875 209.690 ;
        RECT 115.935 206.705 116.165 212.530 ;
        RECT 115.900 206.005 116.200 206.705 ;
        RECT 115.935 204.530 116.165 206.005 ;
        RECT 113.635 203.995 114.595 204.325 ;
        RECT 114.925 203.995 115.885 204.325 ;
        RECT 116.575 203.720 116.975 213.340 ;
        RECT 117.665 212.735 118.625 212.965 ;
        RECT 118.955 212.735 119.915 212.965 ;
        RECT 117.385 205.495 117.615 212.530 ;
        RECT 118.675 211.190 118.905 212.530 ;
        RECT 118.640 209.690 118.940 211.190 ;
        RECT 117.350 204.795 117.650 205.495 ;
        RECT 117.385 204.530 117.615 204.795 ;
        RECT 118.675 204.530 118.905 209.690 ;
        RECT 119.965 206.705 120.195 212.530 ;
        RECT 119.930 206.005 120.230 206.705 ;
        RECT 119.965 204.530 120.195 206.005 ;
        RECT 117.665 203.995 118.625 204.325 ;
        RECT 118.955 203.995 119.915 204.325 ;
        RECT 120.605 203.720 121.005 213.340 ;
        RECT 121.695 212.735 122.655 212.965 ;
        RECT 122.985 212.735 123.945 212.965 ;
        RECT 121.415 205.495 121.645 212.530 ;
        RECT 122.705 211.190 122.935 212.530 ;
        RECT 122.670 209.690 122.970 211.190 ;
        RECT 121.380 204.795 121.680 205.495 ;
        RECT 121.415 204.530 121.645 204.795 ;
        RECT 122.705 204.530 122.935 209.690 ;
        RECT 123.995 206.705 124.225 212.530 ;
        RECT 123.960 206.005 124.260 206.705 ;
        RECT 123.995 204.530 124.225 206.005 ;
        RECT 121.695 203.995 122.655 204.325 ;
        RECT 122.985 203.995 123.945 204.325 ;
        RECT 124.635 203.720 125.035 213.340 ;
        RECT 125.725 212.735 126.685 212.965 ;
        RECT 127.015 212.735 127.975 212.965 ;
        RECT 125.445 205.495 125.675 212.530 ;
        RECT 126.735 211.190 126.965 212.530 ;
        RECT 126.700 209.690 127.000 211.190 ;
        RECT 125.410 204.795 125.710 205.495 ;
        RECT 125.445 204.530 125.675 204.795 ;
        RECT 126.735 204.530 126.965 209.690 ;
        RECT 128.025 206.705 128.255 212.530 ;
        RECT 127.990 206.005 128.290 206.705 ;
        RECT 128.025 204.530 128.255 206.005 ;
        RECT 125.725 203.995 126.685 204.325 ;
        RECT 127.015 203.995 127.975 204.325 ;
        RECT 128.665 203.720 129.065 213.340 ;
        RECT 129.755 212.735 130.715 212.965 ;
        RECT 131.045 212.735 132.005 212.965 ;
        RECT 129.475 205.495 129.705 212.530 ;
        RECT 130.765 211.190 130.995 212.530 ;
        RECT 130.730 209.690 131.030 211.190 ;
        RECT 129.440 204.795 129.740 205.495 ;
        RECT 129.475 204.530 129.705 204.795 ;
        RECT 130.765 204.530 130.995 209.690 ;
        RECT 132.055 206.705 132.285 212.530 ;
        RECT 132.020 206.005 132.320 206.705 ;
        RECT 132.055 204.530 132.285 206.005 ;
        RECT 129.755 203.995 130.715 204.325 ;
        RECT 131.045 203.995 132.005 204.325 ;
        RECT 132.695 203.720 133.095 213.340 ;
        RECT 133.785 212.735 134.745 212.965 ;
        RECT 135.075 212.735 136.035 212.965 ;
        RECT 133.505 205.495 133.735 212.530 ;
        RECT 134.795 211.190 135.025 212.530 ;
        RECT 134.760 209.690 135.060 211.190 ;
        RECT 133.470 204.795 133.770 205.495 ;
        RECT 133.505 204.530 133.735 204.795 ;
        RECT 134.795 204.530 135.025 209.690 ;
        RECT 136.085 206.705 136.315 212.530 ;
        RECT 136.050 206.005 136.350 206.705 ;
        RECT 136.085 204.530 136.315 206.005 ;
        RECT 133.785 203.995 134.745 204.325 ;
        RECT 135.075 203.995 136.035 204.325 ;
        RECT 136.725 203.720 137.125 213.340 ;
        RECT 137.815 212.735 138.775 212.965 ;
        RECT 139.105 212.735 140.065 212.965 ;
        RECT 137.535 205.495 137.765 212.530 ;
        RECT 138.825 211.190 139.055 212.530 ;
        RECT 138.790 209.690 139.090 211.190 ;
        RECT 137.500 204.795 137.800 205.495 ;
        RECT 137.535 204.530 137.765 204.795 ;
        RECT 138.825 204.530 139.055 209.690 ;
        RECT 140.115 206.705 140.345 212.530 ;
        RECT 140.080 206.005 140.380 206.705 ;
        RECT 140.115 204.530 140.345 206.005 ;
        RECT 137.815 203.995 138.775 204.325 ;
        RECT 139.105 203.995 140.065 204.325 ;
        RECT 140.755 203.720 141.155 213.340 ;
        RECT 141.845 212.735 142.805 212.965 ;
        RECT 143.135 212.735 144.095 212.965 ;
        RECT 141.565 205.495 141.795 212.530 ;
        RECT 142.855 211.190 143.085 212.530 ;
        RECT 142.820 209.690 143.120 211.190 ;
        RECT 141.530 204.795 141.830 205.495 ;
        RECT 141.565 204.530 141.795 204.795 ;
        RECT 142.855 204.530 143.085 209.690 ;
        RECT 144.145 206.705 144.375 212.530 ;
        RECT 144.110 206.005 144.410 206.705 ;
        RECT 144.145 204.530 144.375 206.005 ;
        RECT 141.845 203.995 142.805 204.325 ;
        RECT 143.135 203.995 144.095 204.325 ;
        RECT 144.785 203.720 145.185 213.340 ;
        RECT 145.875 212.735 146.835 212.965 ;
        RECT 147.165 212.735 148.125 212.965 ;
        RECT 145.595 205.495 145.825 212.530 ;
        RECT 146.885 211.190 147.115 212.530 ;
        RECT 146.850 209.690 147.150 211.190 ;
        RECT 145.560 204.795 145.860 205.495 ;
        RECT 145.595 204.530 145.825 204.795 ;
        RECT 146.885 204.530 147.115 209.690 ;
        RECT 148.175 206.705 148.405 212.530 ;
        RECT 148.140 206.005 148.440 206.705 ;
        RECT 148.175 204.530 148.405 206.005 ;
        RECT 145.875 203.995 146.835 204.325 ;
        RECT 147.165 203.995 148.125 204.325 ;
        RECT 148.815 203.720 149.215 213.340 ;
        RECT 149.905 212.735 150.865 212.965 ;
        RECT 151.195 212.735 152.155 212.965 ;
        RECT 149.625 205.495 149.855 212.530 ;
        RECT 150.915 211.190 151.145 212.530 ;
        RECT 150.880 209.690 151.180 211.190 ;
        RECT 149.590 204.795 149.890 205.495 ;
        RECT 149.625 204.530 149.855 204.795 ;
        RECT 150.915 204.530 151.145 209.690 ;
        RECT 152.205 206.705 152.435 212.530 ;
        RECT 152.170 206.005 152.470 206.705 ;
        RECT 152.205 204.530 152.435 206.005 ;
        RECT 149.905 203.995 150.865 204.325 ;
        RECT 151.195 203.995 152.155 204.325 ;
        RECT 152.845 203.720 153.245 213.340 ;
        RECT 108.515 203.320 153.245 203.720 ;
        RECT 165.150 201.250 239.210 201.730 ;
        RECT 168.440 201.050 168.760 201.110 ;
        RECT 169.375 201.050 169.665 201.095 ;
        RECT 108.515 200.625 153.245 201.025 ;
        RECT 168.440 200.910 169.665 201.050 ;
        RECT 168.440 200.850 168.760 200.910 ;
        RECT 169.375 200.865 169.665 200.910 ;
        RECT 178.100 201.050 178.420 201.110 ;
        RECT 179.495 201.050 179.785 201.095 ;
        RECT 178.100 200.910 179.785 201.050 ;
        RECT 178.100 200.850 178.420 200.910 ;
        RECT 179.495 200.865 179.785 200.910 ;
        RECT 187.760 201.050 188.080 201.110 ;
        RECT 188.695 201.050 188.985 201.095 ;
        RECT 187.760 200.910 188.985 201.050 ;
        RECT 187.760 200.850 188.080 200.910 ;
        RECT 188.695 200.865 188.985 200.910 ;
        RECT 197.420 201.050 197.740 201.110 ;
        RECT 198.815 201.050 199.105 201.095 ;
        RECT 197.420 200.910 199.105 201.050 ;
        RECT 197.420 200.850 197.740 200.910 ;
        RECT 198.815 200.865 199.105 200.910 ;
        RECT 207.080 201.050 207.400 201.110 ;
        RECT 208.015 201.050 208.305 201.095 ;
        RECT 207.080 200.910 208.305 201.050 ;
        RECT 207.080 200.850 207.400 200.910 ;
        RECT 208.015 200.865 208.305 200.910 ;
        RECT 216.740 201.050 217.060 201.110 ;
        RECT 218.135 201.050 218.425 201.095 ;
        RECT 216.740 200.910 218.425 201.050 ;
        RECT 216.740 200.850 217.060 200.910 ;
        RECT 218.135 200.865 218.425 200.910 ;
        RECT 226.400 201.050 226.720 201.110 ;
        RECT 227.795 201.050 228.085 201.095 ;
        RECT 226.400 200.910 228.085 201.050 ;
        RECT 226.400 200.850 226.720 200.910 ;
        RECT 227.795 200.865 228.085 200.910 ;
        RECT 236.060 201.050 236.380 201.110 ;
        RECT 236.995 201.050 237.285 201.095 ;
        RECT 236.060 200.910 237.285 201.050 ;
        RECT 236.060 200.850 236.380 200.910 ;
        RECT 236.995 200.865 237.285 200.910 ;
        RECT 108.515 195.095 108.915 200.625 ;
        RECT 109.735 200.250 110.435 200.320 ;
        RECT 111.025 200.250 111.725 200.320 ;
        RECT 109.605 200.020 110.565 200.250 ;
        RECT 110.895 200.020 111.855 200.250 ;
        RECT 109.325 199.635 109.555 199.860 ;
        RECT 109.290 198.935 109.590 199.635 ;
        RECT 110.615 198.955 110.845 199.860 ;
        RECT 111.905 199.635 112.135 199.860 ;
        RECT 109.325 195.860 109.555 198.935 ;
        RECT 110.580 196.855 110.880 198.955 ;
        RECT 111.870 198.935 112.170 199.635 ;
        RECT 110.615 195.860 110.845 196.855 ;
        RECT 111.905 195.860 112.135 198.935 ;
        RECT 109.605 195.470 110.565 195.700 ;
        RECT 110.895 195.470 111.855 195.700 ;
        RECT 112.545 195.095 112.945 200.625 ;
        RECT 113.765 200.250 114.465 200.320 ;
        RECT 115.055 200.250 115.755 200.320 ;
        RECT 113.635 200.020 114.595 200.250 ;
        RECT 114.925 200.020 115.885 200.250 ;
        RECT 113.355 199.635 113.585 199.860 ;
        RECT 113.320 198.935 113.620 199.635 ;
        RECT 114.645 198.955 114.875 199.860 ;
        RECT 115.935 199.635 116.165 199.860 ;
        RECT 113.355 195.860 113.585 198.935 ;
        RECT 114.610 196.855 114.910 198.955 ;
        RECT 115.900 198.935 116.200 199.635 ;
        RECT 114.645 195.860 114.875 196.855 ;
        RECT 115.935 195.860 116.165 198.935 ;
        RECT 113.635 195.470 114.595 195.700 ;
        RECT 114.925 195.470 115.885 195.700 ;
        RECT 116.575 195.095 116.975 200.625 ;
        RECT 117.795 200.250 118.495 200.320 ;
        RECT 119.085 200.250 119.785 200.320 ;
        RECT 117.665 200.020 118.625 200.250 ;
        RECT 118.955 200.020 119.915 200.250 ;
        RECT 117.385 199.635 117.615 199.860 ;
        RECT 117.350 198.935 117.650 199.635 ;
        RECT 118.675 198.955 118.905 199.860 ;
        RECT 119.965 199.635 120.195 199.860 ;
        RECT 117.385 195.860 117.615 198.935 ;
        RECT 118.640 196.855 118.940 198.955 ;
        RECT 119.930 198.935 120.230 199.635 ;
        RECT 118.675 195.860 118.905 196.855 ;
        RECT 119.965 195.860 120.195 198.935 ;
        RECT 117.665 195.470 118.625 195.700 ;
        RECT 118.955 195.470 119.915 195.700 ;
        RECT 120.605 195.095 121.005 200.625 ;
        RECT 121.825 200.250 122.525 200.320 ;
        RECT 123.115 200.250 123.815 200.320 ;
        RECT 121.695 200.020 122.655 200.250 ;
        RECT 122.985 200.020 123.945 200.250 ;
        RECT 121.415 199.635 121.645 199.860 ;
        RECT 121.380 198.935 121.680 199.635 ;
        RECT 122.705 198.955 122.935 199.860 ;
        RECT 123.995 199.635 124.225 199.860 ;
        RECT 121.415 195.860 121.645 198.935 ;
        RECT 122.670 196.855 122.970 198.955 ;
        RECT 123.960 198.935 124.260 199.635 ;
        RECT 122.705 195.860 122.935 196.855 ;
        RECT 123.995 195.860 124.225 198.935 ;
        RECT 121.695 195.470 122.655 195.700 ;
        RECT 122.985 195.470 123.945 195.700 ;
        RECT 124.635 195.095 125.035 200.625 ;
        RECT 125.855 200.250 126.555 200.320 ;
        RECT 127.145 200.250 127.845 200.320 ;
        RECT 125.725 200.020 126.685 200.250 ;
        RECT 127.015 200.020 127.975 200.250 ;
        RECT 125.445 199.635 125.675 199.860 ;
        RECT 125.410 198.935 125.710 199.635 ;
        RECT 126.735 198.955 126.965 199.860 ;
        RECT 128.025 199.635 128.255 199.860 ;
        RECT 125.445 195.860 125.675 198.935 ;
        RECT 126.700 196.855 127.000 198.955 ;
        RECT 127.990 198.935 128.290 199.635 ;
        RECT 126.735 195.860 126.965 196.855 ;
        RECT 128.025 195.860 128.255 198.935 ;
        RECT 125.725 195.470 126.685 195.700 ;
        RECT 127.015 195.470 127.975 195.700 ;
        RECT 128.665 195.095 129.065 200.625 ;
        RECT 129.885 200.250 130.585 200.320 ;
        RECT 131.175 200.250 131.875 200.320 ;
        RECT 129.755 200.020 130.715 200.250 ;
        RECT 131.045 200.020 132.005 200.250 ;
        RECT 129.475 199.635 129.705 199.860 ;
        RECT 129.440 198.935 129.740 199.635 ;
        RECT 130.765 198.955 130.995 199.860 ;
        RECT 132.055 199.635 132.285 199.860 ;
        RECT 129.475 195.860 129.705 198.935 ;
        RECT 130.730 196.855 131.030 198.955 ;
        RECT 132.020 198.935 132.320 199.635 ;
        RECT 130.765 195.860 130.995 196.855 ;
        RECT 132.055 195.860 132.285 198.935 ;
        RECT 129.755 195.470 130.715 195.700 ;
        RECT 131.045 195.470 132.005 195.700 ;
        RECT 132.695 195.095 133.095 200.625 ;
        RECT 133.915 200.250 134.615 200.320 ;
        RECT 135.205 200.250 135.905 200.320 ;
        RECT 133.785 200.020 134.745 200.250 ;
        RECT 135.075 200.020 136.035 200.250 ;
        RECT 133.505 199.635 133.735 199.860 ;
        RECT 133.470 198.935 133.770 199.635 ;
        RECT 134.795 198.955 135.025 199.860 ;
        RECT 136.085 199.635 136.315 199.860 ;
        RECT 133.505 195.860 133.735 198.935 ;
        RECT 134.760 196.855 135.060 198.955 ;
        RECT 136.050 198.935 136.350 199.635 ;
        RECT 134.795 195.860 135.025 196.855 ;
        RECT 136.085 195.860 136.315 198.935 ;
        RECT 133.785 195.470 134.745 195.700 ;
        RECT 135.075 195.470 136.035 195.700 ;
        RECT 136.725 195.095 137.125 200.625 ;
        RECT 137.945 200.250 138.645 200.320 ;
        RECT 139.235 200.250 139.935 200.320 ;
        RECT 137.815 200.020 138.775 200.250 ;
        RECT 139.105 200.020 140.065 200.250 ;
        RECT 137.535 199.635 137.765 199.860 ;
        RECT 137.500 198.935 137.800 199.635 ;
        RECT 138.825 198.955 139.055 199.860 ;
        RECT 140.115 199.635 140.345 199.860 ;
        RECT 137.535 195.860 137.765 198.935 ;
        RECT 138.790 196.855 139.090 198.955 ;
        RECT 140.080 198.935 140.380 199.635 ;
        RECT 138.825 195.860 139.055 196.855 ;
        RECT 140.115 195.860 140.345 198.935 ;
        RECT 137.815 195.470 138.775 195.700 ;
        RECT 139.105 195.470 140.065 195.700 ;
        RECT 140.755 195.095 141.155 200.625 ;
        RECT 141.975 200.250 142.675 200.320 ;
        RECT 143.265 200.250 143.965 200.320 ;
        RECT 141.845 200.020 142.805 200.250 ;
        RECT 143.135 200.020 144.095 200.250 ;
        RECT 141.565 199.635 141.795 199.860 ;
        RECT 141.530 198.935 141.830 199.635 ;
        RECT 142.855 198.955 143.085 199.860 ;
        RECT 144.145 199.635 144.375 199.860 ;
        RECT 141.565 195.860 141.795 198.935 ;
        RECT 142.820 196.855 143.120 198.955 ;
        RECT 144.110 198.935 144.410 199.635 ;
        RECT 142.855 195.860 143.085 196.855 ;
        RECT 144.145 195.860 144.375 198.935 ;
        RECT 141.845 195.470 142.805 195.700 ;
        RECT 143.135 195.470 144.095 195.700 ;
        RECT 144.785 195.095 145.185 200.625 ;
        RECT 146.005 200.250 146.705 200.320 ;
        RECT 147.295 200.250 147.995 200.320 ;
        RECT 145.875 200.020 146.835 200.250 ;
        RECT 147.165 200.020 148.125 200.250 ;
        RECT 145.595 199.635 145.825 199.860 ;
        RECT 145.560 198.935 145.860 199.635 ;
        RECT 146.885 198.955 147.115 199.860 ;
        RECT 148.175 199.635 148.405 199.860 ;
        RECT 145.595 195.860 145.825 198.935 ;
        RECT 146.850 196.855 147.150 198.955 ;
        RECT 148.140 198.935 148.440 199.635 ;
        RECT 146.885 195.860 147.115 196.855 ;
        RECT 148.175 195.860 148.405 198.935 ;
        RECT 145.875 195.470 146.835 195.700 ;
        RECT 147.165 195.470 148.125 195.700 ;
        RECT 148.815 195.095 149.215 200.625 ;
        RECT 150.035 200.250 150.735 200.320 ;
        RECT 151.325 200.250 152.025 200.320 ;
        RECT 149.905 200.020 150.865 200.250 ;
        RECT 151.195 200.020 152.155 200.250 ;
        RECT 149.625 199.635 149.855 199.860 ;
        RECT 149.590 198.935 149.890 199.635 ;
        RECT 150.915 198.955 151.145 199.860 ;
        RECT 152.205 199.635 152.435 199.860 ;
        RECT 149.625 195.860 149.855 198.935 ;
        RECT 150.880 196.855 151.180 198.955 ;
        RECT 152.170 198.935 152.470 199.635 ;
        RECT 150.915 195.860 151.145 196.855 ;
        RECT 152.205 195.860 152.435 198.935 ;
        RECT 149.905 195.470 150.865 195.700 ;
        RECT 151.195 195.470 152.155 195.700 ;
        RECT 152.845 195.095 153.245 200.625 ;
        RECT 166.600 199.830 166.920 200.090 ;
        RECT 170.280 199.830 170.600 200.090 ;
        RECT 178.560 199.830 178.880 200.090 ;
        RECT 189.615 200.030 189.905 200.075 ;
        RECT 191.440 200.030 191.760 200.090 ;
        RECT 189.615 199.890 191.760 200.030 ;
        RECT 189.615 199.845 189.905 199.890 ;
        RECT 191.440 199.830 191.760 199.890 ;
        RECT 197.880 199.830 198.200 200.090 ;
        RECT 208.920 199.830 209.240 200.090 ;
        RECT 217.200 199.830 217.520 200.090 ;
        RECT 226.860 199.830 227.180 200.090 ;
        RECT 236.060 199.830 236.380 200.090 ;
        RECT 167.535 199.350 167.825 199.395 ;
        RECT 174.420 199.350 174.740 199.410 ;
        RECT 167.535 199.210 174.740 199.350 ;
        RECT 167.535 199.165 167.825 199.210 ;
        RECT 174.420 199.150 174.740 199.210 ;
        RECT 165.150 198.530 239.210 199.010 ;
        RECT 165.150 195.810 239.210 196.290 ;
        RECT 108.515 194.695 153.245 195.095 ;
        RECT 108.515 185.165 108.915 194.695 ;
        RECT 109.605 194.320 110.305 194.390 ;
        RECT 111.155 194.320 111.855 194.390 ;
        RECT 109.605 194.090 110.565 194.320 ;
        RECT 110.895 194.090 111.855 194.320 ;
        RECT 109.325 192.835 109.555 193.930 ;
        RECT 109.290 191.335 109.590 192.835 ;
        RECT 109.325 185.930 109.555 191.335 ;
        RECT 110.615 189.090 110.845 193.930 ;
        RECT 111.905 192.835 112.135 193.930 ;
        RECT 111.870 191.335 112.170 192.835 ;
        RECT 110.580 187.590 110.880 189.090 ;
        RECT 110.615 185.930 110.845 187.590 ;
        RECT 111.905 185.930 112.135 191.335 ;
        RECT 109.605 185.540 110.565 185.770 ;
        RECT 110.895 185.540 111.855 185.770 ;
        RECT 112.545 185.165 112.945 194.695 ;
        RECT 113.635 194.320 114.335 194.390 ;
        RECT 115.185 194.320 115.885 194.390 ;
        RECT 113.635 194.090 114.595 194.320 ;
        RECT 114.925 194.090 115.885 194.320 ;
        RECT 113.355 192.835 113.585 193.930 ;
        RECT 113.320 191.335 113.620 192.835 ;
        RECT 113.355 185.930 113.585 191.335 ;
        RECT 114.645 189.090 114.875 193.930 ;
        RECT 115.935 192.835 116.165 193.930 ;
        RECT 115.900 191.335 116.200 192.835 ;
        RECT 114.610 187.590 114.910 189.090 ;
        RECT 114.645 185.930 114.875 187.590 ;
        RECT 115.935 185.930 116.165 191.335 ;
        RECT 113.635 185.540 114.595 185.770 ;
        RECT 114.925 185.540 115.885 185.770 ;
        RECT 116.575 185.165 116.975 194.695 ;
        RECT 117.665 194.320 118.365 194.390 ;
        RECT 119.215 194.320 119.915 194.390 ;
        RECT 117.665 194.090 118.625 194.320 ;
        RECT 118.955 194.090 119.915 194.320 ;
        RECT 117.385 192.835 117.615 193.930 ;
        RECT 117.350 191.335 117.650 192.835 ;
        RECT 117.385 185.930 117.615 191.335 ;
        RECT 118.675 189.090 118.905 193.930 ;
        RECT 119.965 192.835 120.195 193.930 ;
        RECT 119.930 191.335 120.230 192.835 ;
        RECT 118.640 187.590 118.940 189.090 ;
        RECT 118.675 185.930 118.905 187.590 ;
        RECT 119.965 185.930 120.195 191.335 ;
        RECT 117.665 185.540 118.625 185.770 ;
        RECT 118.955 185.540 119.915 185.770 ;
        RECT 120.605 185.165 121.005 194.695 ;
        RECT 121.695 194.320 122.395 194.390 ;
        RECT 123.245 194.320 123.945 194.390 ;
        RECT 121.695 194.090 122.655 194.320 ;
        RECT 122.985 194.090 123.945 194.320 ;
        RECT 121.415 192.835 121.645 193.930 ;
        RECT 121.380 191.335 121.680 192.835 ;
        RECT 121.415 185.930 121.645 191.335 ;
        RECT 122.705 189.090 122.935 193.930 ;
        RECT 123.995 192.835 124.225 193.930 ;
        RECT 123.960 191.335 124.260 192.835 ;
        RECT 122.670 187.590 122.970 189.090 ;
        RECT 122.705 185.930 122.935 187.590 ;
        RECT 123.995 185.930 124.225 191.335 ;
        RECT 121.695 185.540 122.655 185.770 ;
        RECT 122.985 185.540 123.945 185.770 ;
        RECT 124.635 185.165 125.035 194.695 ;
        RECT 125.725 194.320 126.425 194.390 ;
        RECT 127.275 194.320 127.975 194.390 ;
        RECT 125.725 194.090 126.685 194.320 ;
        RECT 127.015 194.090 127.975 194.320 ;
        RECT 125.445 192.835 125.675 193.930 ;
        RECT 125.410 191.335 125.710 192.835 ;
        RECT 125.445 185.930 125.675 191.335 ;
        RECT 126.735 189.090 126.965 193.930 ;
        RECT 128.025 192.835 128.255 193.930 ;
        RECT 127.990 191.335 128.290 192.835 ;
        RECT 126.700 187.590 127.000 189.090 ;
        RECT 126.735 185.930 126.965 187.590 ;
        RECT 128.025 185.930 128.255 191.335 ;
        RECT 125.725 185.540 126.685 185.770 ;
        RECT 127.015 185.540 127.975 185.770 ;
        RECT 128.665 185.165 129.065 194.695 ;
        RECT 129.755 194.320 130.455 194.390 ;
        RECT 131.305 194.320 132.005 194.390 ;
        RECT 129.755 194.090 130.715 194.320 ;
        RECT 131.045 194.090 132.005 194.320 ;
        RECT 129.475 192.835 129.705 193.930 ;
        RECT 129.440 191.335 129.740 192.835 ;
        RECT 129.475 185.930 129.705 191.335 ;
        RECT 130.765 189.090 130.995 193.930 ;
        RECT 132.055 192.835 132.285 193.930 ;
        RECT 132.020 191.335 132.320 192.835 ;
        RECT 130.730 187.590 131.030 189.090 ;
        RECT 130.765 185.930 130.995 187.590 ;
        RECT 132.055 185.930 132.285 191.335 ;
        RECT 129.755 185.540 130.715 185.770 ;
        RECT 131.045 185.540 132.005 185.770 ;
        RECT 132.695 185.165 133.095 194.695 ;
        RECT 133.785 194.320 134.485 194.390 ;
        RECT 135.335 194.320 136.035 194.390 ;
        RECT 133.785 194.090 134.745 194.320 ;
        RECT 135.075 194.090 136.035 194.320 ;
        RECT 133.505 192.835 133.735 193.930 ;
        RECT 133.470 191.335 133.770 192.835 ;
        RECT 133.505 185.930 133.735 191.335 ;
        RECT 134.795 189.090 135.025 193.930 ;
        RECT 136.085 192.835 136.315 193.930 ;
        RECT 136.050 191.335 136.350 192.835 ;
        RECT 134.760 187.590 135.060 189.090 ;
        RECT 134.795 185.930 135.025 187.590 ;
        RECT 136.085 185.930 136.315 191.335 ;
        RECT 133.785 185.540 134.745 185.770 ;
        RECT 135.075 185.540 136.035 185.770 ;
        RECT 136.725 185.165 137.125 194.695 ;
        RECT 137.815 194.320 138.515 194.390 ;
        RECT 139.365 194.320 140.065 194.390 ;
        RECT 137.815 194.090 138.775 194.320 ;
        RECT 139.105 194.090 140.065 194.320 ;
        RECT 137.535 192.835 137.765 193.930 ;
        RECT 137.500 191.335 137.800 192.835 ;
        RECT 137.535 185.930 137.765 191.335 ;
        RECT 138.825 189.090 139.055 193.930 ;
        RECT 140.115 192.835 140.345 193.930 ;
        RECT 140.080 191.335 140.380 192.835 ;
        RECT 138.790 187.590 139.090 189.090 ;
        RECT 138.825 185.930 139.055 187.590 ;
        RECT 140.115 185.930 140.345 191.335 ;
        RECT 137.815 185.540 138.775 185.770 ;
        RECT 139.105 185.540 140.065 185.770 ;
        RECT 140.755 185.165 141.155 194.695 ;
        RECT 141.845 194.320 142.545 194.390 ;
        RECT 143.395 194.320 144.095 194.390 ;
        RECT 141.845 194.090 142.805 194.320 ;
        RECT 143.135 194.090 144.095 194.320 ;
        RECT 141.565 192.835 141.795 193.930 ;
        RECT 141.530 191.335 141.830 192.835 ;
        RECT 141.565 185.930 141.795 191.335 ;
        RECT 142.855 189.090 143.085 193.930 ;
        RECT 144.145 192.835 144.375 193.930 ;
        RECT 144.110 191.335 144.410 192.835 ;
        RECT 142.820 187.590 143.120 189.090 ;
        RECT 142.855 185.930 143.085 187.590 ;
        RECT 144.145 185.930 144.375 191.335 ;
        RECT 141.845 185.540 142.805 185.770 ;
        RECT 143.135 185.540 144.095 185.770 ;
        RECT 144.785 185.165 145.185 194.695 ;
        RECT 145.875 194.320 146.575 194.390 ;
        RECT 147.425 194.320 148.125 194.390 ;
        RECT 145.875 194.090 146.835 194.320 ;
        RECT 147.165 194.090 148.125 194.320 ;
        RECT 145.595 192.835 145.825 193.930 ;
        RECT 145.560 191.335 145.860 192.835 ;
        RECT 145.595 185.930 145.825 191.335 ;
        RECT 146.885 189.090 147.115 193.930 ;
        RECT 148.175 192.835 148.405 193.930 ;
        RECT 148.140 191.335 148.440 192.835 ;
        RECT 146.850 187.590 147.150 189.090 ;
        RECT 146.885 185.930 147.115 187.590 ;
        RECT 148.175 185.930 148.405 191.335 ;
        RECT 145.875 185.540 146.835 185.770 ;
        RECT 147.165 185.540 148.125 185.770 ;
        RECT 148.815 185.165 149.215 194.695 ;
        RECT 149.905 194.320 150.605 194.390 ;
        RECT 151.455 194.320 152.155 194.390 ;
        RECT 149.905 194.090 150.865 194.320 ;
        RECT 151.195 194.090 152.155 194.320 ;
        RECT 149.625 192.835 149.855 193.930 ;
        RECT 149.590 191.335 149.890 192.835 ;
        RECT 149.625 185.930 149.855 191.335 ;
        RECT 150.915 189.090 151.145 193.930 ;
        RECT 152.205 192.835 152.435 193.930 ;
        RECT 152.170 191.335 152.470 192.835 ;
        RECT 150.880 187.590 151.180 189.090 ;
        RECT 150.915 185.930 151.145 187.590 ;
        RECT 152.205 185.930 152.435 191.335 ;
        RECT 152.845 187.965 153.245 194.695 ;
        RECT 181.320 193.910 181.640 193.970 ;
        RECT 207.540 193.910 207.860 193.970 ;
        RECT 181.320 193.770 207.860 193.910 ;
        RECT 181.320 193.710 181.640 193.770 ;
        RECT 207.540 193.710 207.860 193.770 ;
        RECT 165.150 193.090 239.210 193.570 ;
        RECT 177.655 192.890 177.945 192.935 ;
        RECT 178.560 192.890 178.880 192.950 ;
        RECT 177.655 192.750 178.880 192.890 ;
        RECT 177.655 192.705 177.945 192.750 ;
        RECT 178.560 192.690 178.880 192.750 ;
        RECT 182.240 192.890 182.560 192.950 ;
        RECT 182.240 192.750 188.910 192.890 ;
        RECT 182.240 192.690 182.560 192.750 ;
        RECT 181.780 192.550 182.100 192.610 ;
        RECT 180.490 192.410 182.100 192.550 ;
        RECT 173.500 192.210 173.820 192.270 ;
        RECT 173.975 192.210 174.265 192.255 ;
        RECT 173.500 192.070 174.265 192.210 ;
        RECT 173.500 192.010 173.820 192.070 ;
        RECT 173.975 192.025 174.265 192.070 ;
        RECT 174.435 192.210 174.725 192.255 ;
        RECT 175.340 192.210 175.660 192.270 ;
        RECT 174.435 192.070 175.660 192.210 ;
        RECT 174.435 192.025 174.725 192.070 ;
        RECT 175.340 192.010 175.660 192.070 ;
        RECT 176.735 192.210 177.025 192.255 ;
        RECT 177.640 192.210 177.960 192.270 ;
        RECT 176.735 192.070 177.960 192.210 ;
        RECT 176.735 192.025 177.025 192.070 ;
        RECT 177.640 192.010 177.960 192.070 ;
        RECT 178.560 192.010 178.880 192.270 ;
        RECT 179.020 192.200 179.340 192.270 ;
        RECT 180.490 192.255 180.630 192.410 ;
        RECT 181.780 192.350 182.100 192.410 ;
        RECT 185.475 192.550 185.765 192.595 ;
        RECT 188.220 192.550 188.540 192.610 ;
        RECT 185.475 192.410 188.540 192.550 ;
        RECT 188.770 192.550 188.910 192.750 ;
        RECT 191.440 192.690 191.760 192.950 ;
        RECT 197.880 192.690 198.200 192.950 ;
        RECT 216.740 192.550 217.060 192.610 ;
        RECT 188.770 192.410 217.060 192.550 ;
        RECT 185.475 192.365 185.765 192.410 ;
        RECT 188.220 192.350 188.540 192.410 ;
        RECT 216.740 192.350 217.060 192.410 ;
        RECT 179.935 192.210 180.225 192.255 ;
        RECT 179.805 192.200 180.225 192.210 ;
        RECT 179.020 192.060 180.225 192.200 ;
        RECT 179.020 192.010 179.340 192.060 ;
        RECT 179.935 192.025 180.225 192.060 ;
        RECT 180.415 192.025 180.705 192.255 ;
        RECT 180.860 192.210 181.180 192.270 ;
        RECT 182.255 192.210 182.545 192.255 ;
        RECT 180.860 192.070 182.545 192.210 ;
        RECT 180.860 192.010 181.180 192.070 ;
        RECT 182.255 192.025 182.545 192.070 ;
        RECT 184.080 192.010 184.400 192.270 ;
        RECT 184.560 192.025 184.850 192.255 ;
        RECT 179.495 191.870 179.785 191.915 ;
        RECT 181.780 191.870 182.100 191.930 ;
        RECT 179.495 191.730 182.100 191.870 ;
        RECT 179.495 191.685 179.785 191.730 ;
        RECT 181.780 191.670 182.100 191.730 ;
        RECT 182.700 191.870 183.020 191.930 ;
        RECT 184.635 191.870 184.775 192.025 ;
        RECT 185.920 192.010 186.240 192.270 ;
        RECT 186.420 192.025 186.710 192.255 ;
        RECT 192.375 192.210 192.665 192.255 ;
        RECT 187.390 192.070 192.665 192.210 ;
        RECT 182.700 191.730 184.775 191.870 ;
        RECT 182.700 191.670 183.020 191.730 ;
        RECT 175.800 191.330 176.120 191.590 ;
        RECT 178.100 191.530 178.420 191.590 ;
        RECT 186.470 191.530 186.610 192.025 ;
        RECT 187.390 191.575 187.530 192.070 ;
        RECT 192.375 192.025 192.665 192.070 ;
        RECT 194.200 192.210 194.520 192.270 ;
        RECT 197.435 192.210 197.725 192.255 ;
        RECT 194.200 192.070 197.725 192.210 ;
        RECT 194.200 192.010 194.520 192.070 ;
        RECT 197.435 192.025 197.725 192.070 ;
        RECT 198.800 192.010 199.120 192.270 ;
        RECT 193.740 191.870 194.060 191.930 ;
        RECT 196.975 191.870 197.265 191.915 ;
        RECT 200.180 191.870 200.500 191.930 ;
        RECT 193.740 191.730 200.500 191.870 ;
        RECT 193.740 191.670 194.060 191.730 ;
        RECT 196.975 191.685 197.265 191.730 ;
        RECT 200.180 191.670 200.500 191.730 ;
        RECT 178.100 191.390 186.610 191.530 ;
        RECT 178.100 191.330 178.420 191.390 ;
        RECT 187.315 191.345 187.605 191.575 ;
        RECT 193.295 191.530 193.585 191.575 ;
        RECT 206.620 191.530 206.940 191.590 ;
        RECT 193.295 191.390 206.940 191.530 ;
        RECT 193.295 191.345 193.585 191.390 ;
        RECT 206.620 191.330 206.940 191.390 ;
        RECT 173.040 190.990 173.360 191.250 ;
        RECT 174.880 191.190 175.200 191.250 ;
        RECT 175.355 191.190 175.645 191.235 ;
        RECT 174.880 191.050 175.645 191.190 ;
        RECT 174.880 190.990 175.200 191.050 ;
        RECT 175.355 191.005 175.645 191.050 ;
        RECT 177.640 191.190 177.960 191.250 ;
        RECT 181.320 191.190 181.640 191.250 ;
        RECT 177.640 191.050 181.640 191.190 ;
        RECT 177.640 190.990 177.960 191.050 ;
        RECT 181.320 190.990 181.640 191.050 ;
        RECT 183.160 190.990 183.480 191.250 ;
        RECT 199.735 191.190 200.025 191.235 ;
        RECT 202.940 191.190 203.260 191.250 ;
        RECT 199.735 191.050 203.260 191.190 ;
        RECT 199.735 191.005 200.025 191.050 ;
        RECT 202.940 190.990 203.260 191.050 ;
        RECT 225.940 191.190 226.260 191.250 ;
        RECT 232.380 191.190 232.700 191.250 ;
        RECT 225.940 191.050 232.700 191.190 ;
        RECT 225.940 190.990 226.260 191.050 ;
        RECT 232.380 190.990 232.700 191.050 ;
        RECT 165.150 190.370 239.210 190.850 ;
        RECT 167.520 189.970 167.840 190.230 ;
        RECT 170.280 190.170 170.600 190.230 ;
        RECT 171.215 190.170 171.505 190.215 ;
        RECT 170.280 190.030 171.505 190.170 ;
        RECT 170.280 189.970 170.600 190.030 ;
        RECT 171.215 189.985 171.505 190.030 ;
        RECT 181.795 190.170 182.085 190.215 ;
        RECT 192.835 190.170 193.125 190.215 ;
        RECT 198.800 190.170 199.120 190.230 ;
        RECT 181.795 190.030 188.910 190.170 ;
        RECT 181.795 189.985 182.085 190.030 ;
        RECT 173.960 189.830 174.280 189.890 ;
        RECT 169.910 189.690 174.280 189.830 ;
        RECT 166.600 188.950 166.920 189.210 ;
        RECT 169.910 189.195 170.050 189.690 ;
        RECT 173.960 189.630 174.280 189.690 ;
        RECT 184.555 189.830 184.845 189.875 ;
        RECT 185.920 189.830 186.240 189.890 ;
        RECT 184.555 189.690 186.240 189.830 ;
        RECT 184.555 189.645 184.845 189.690 ;
        RECT 185.920 189.630 186.240 189.690 ;
        RECT 171.660 189.490 171.980 189.550 ;
        RECT 173.055 189.490 173.345 189.535 ;
        RECT 171.660 189.350 173.345 189.490 ;
        RECT 171.660 189.290 171.980 189.350 ;
        RECT 173.055 189.305 173.345 189.350 ;
        RECT 173.515 189.490 173.805 189.535 ;
        RECT 179.020 189.490 179.340 189.550 ;
        RECT 185.000 189.490 185.320 189.550 ;
        RECT 188.770 189.490 188.910 190.030 ;
        RECT 192.835 190.030 199.120 190.170 ;
        RECT 192.835 189.985 193.125 190.030 ;
        RECT 198.800 189.970 199.120 190.030 ;
        RECT 216.295 190.170 216.585 190.215 ;
        RECT 217.200 190.170 217.520 190.230 ;
        RECT 216.295 190.030 217.520 190.170 ;
        RECT 216.295 189.985 216.585 190.030 ;
        RECT 217.200 189.970 217.520 190.030 ;
        RECT 218.135 190.170 218.425 190.215 ;
        RECT 225.940 190.170 226.260 190.230 ;
        RECT 218.135 190.030 226.260 190.170 ;
        RECT 218.135 189.985 218.425 190.030 ;
        RECT 225.940 189.970 226.260 190.030 ;
        RECT 226.415 190.170 226.705 190.215 ;
        RECT 226.860 190.170 227.180 190.230 ;
        RECT 232.855 190.170 233.145 190.215 ;
        RECT 226.415 190.030 227.180 190.170 ;
        RECT 226.415 189.985 226.705 190.030 ;
        RECT 226.860 189.970 227.180 190.030 ;
        RECT 227.410 190.030 233.145 190.170 ;
        RECT 225.020 189.830 225.340 189.890 ;
        RECT 227.410 189.830 227.550 190.030 ;
        RECT 232.855 189.985 233.145 190.030 ;
        RECT 225.020 189.690 227.550 189.830 ;
        RECT 231.015 189.830 231.305 189.875 ;
        RECT 231.460 189.830 231.780 189.890 ;
        RECT 231.015 189.690 231.780 189.830 ;
        RECT 225.020 189.630 225.340 189.690 ;
        RECT 231.015 189.645 231.305 189.690 ;
        RECT 231.460 189.630 231.780 189.690 ;
        RECT 200.180 189.490 200.500 189.550 ;
        RECT 210.300 189.490 210.620 189.550 ;
        RECT 218.595 189.490 218.885 189.535 ;
        RECT 228.715 189.490 229.005 189.535 ;
        RECT 230.540 189.490 230.860 189.550 ;
        RECT 173.515 189.350 179.340 189.490 ;
        RECT 173.515 189.305 173.805 189.350 ;
        RECT 179.020 189.290 179.340 189.350 ;
        RECT 180.490 189.350 183.395 189.490 ;
        RECT 169.835 188.965 170.125 189.195 ;
        RECT 172.120 188.950 172.440 189.210 ;
        RECT 173.975 188.965 174.265 189.195 ;
        RECT 174.050 188.810 174.190 188.965 ;
        RECT 174.880 188.950 175.200 189.210 ;
        RECT 176.260 188.950 176.580 189.210 ;
        RECT 178.575 188.965 178.865 189.195 ;
        RECT 179.495 189.150 179.785 189.195 ;
        RECT 179.940 189.150 180.260 189.210 ;
        RECT 179.495 189.010 180.260 189.150 ;
        RECT 179.495 188.965 179.785 189.010 ;
        RECT 177.640 188.810 177.960 188.870 ;
        RECT 178.650 188.810 178.790 188.965 ;
        RECT 179.940 188.950 180.260 189.010 ;
        RECT 180.490 188.810 180.630 189.350 ;
        RECT 180.860 189.150 181.180 189.210 ;
        RECT 182.240 189.150 182.560 189.210 ;
        RECT 183.255 189.195 183.395 189.350 ;
        RECT 185.000 189.350 188.450 189.490 ;
        RECT 188.770 189.350 192.155 189.490 ;
        RECT 185.000 189.290 185.320 189.350 ;
        RECT 180.860 189.010 182.560 189.150 ;
        RECT 180.860 188.950 181.180 189.010 ;
        RECT 182.240 188.950 182.560 189.010 ;
        RECT 182.715 188.965 183.005 189.195 ;
        RECT 183.180 188.965 183.470 189.195 ;
        RECT 185.935 188.965 186.225 189.195 ;
        RECT 174.050 188.670 180.630 188.810 ;
        RECT 177.640 188.610 177.960 188.670 ;
        RECT 170.755 188.470 171.045 188.515 ;
        RECT 172.580 188.470 172.900 188.530 ;
        RECT 170.755 188.330 172.900 188.470 ;
        RECT 170.755 188.285 171.045 188.330 ;
        RECT 172.580 188.270 172.900 188.330 ;
        RECT 177.195 188.470 177.485 188.515 ;
        RECT 178.100 188.470 178.420 188.530 ;
        RECT 177.195 188.330 178.420 188.470 ;
        RECT 177.195 188.285 177.485 188.330 ;
        RECT 178.100 188.270 178.420 188.330 ;
        RECT 182.240 188.470 182.560 188.530 ;
        RECT 182.790 188.470 182.930 188.965 ;
        RECT 182.240 188.330 182.930 188.470 ;
        RECT 182.240 188.270 182.560 188.330 ;
        RECT 185.000 188.270 185.320 188.530 ;
        RECT 186.010 188.470 186.150 188.965 ;
        RECT 186.380 188.950 186.700 189.210 ;
        RECT 186.840 189.150 187.160 189.210 ;
        RECT 188.310 189.150 188.450 189.350 ;
        RECT 189.140 189.150 189.460 189.210 ;
        RECT 189.615 189.150 189.905 189.195 ;
        RECT 186.840 189.010 187.355 189.150 ;
        RECT 188.310 189.010 189.905 189.150 ;
        RECT 186.840 188.950 187.160 189.010 ;
        RECT 189.140 188.950 189.460 189.010 ;
        RECT 189.615 188.965 189.905 189.010 ;
        RECT 190.060 189.150 190.380 189.210 ;
        RECT 190.060 189.010 190.575 189.150 ;
        RECT 190.060 188.950 190.380 189.010 ;
        RECT 190.980 188.950 191.300 189.210 ;
        RECT 192.015 189.195 192.155 189.350 ;
        RECT 200.180 189.350 230.860 189.490 ;
        RECT 200.180 189.290 200.500 189.350 ;
        RECT 210.300 189.290 210.620 189.350 ;
        RECT 218.595 189.305 218.885 189.350 ;
        RECT 228.715 189.305 229.005 189.350 ;
        RECT 230.540 189.290 230.860 189.350 ;
        RECT 191.940 188.965 192.230 189.195 ;
        RECT 196.500 188.950 196.820 189.210 ;
        RECT 196.980 188.965 197.270 189.195 ;
        RECT 210.760 189.150 211.080 189.210 ;
        RECT 217.215 189.150 217.505 189.195 ;
        RECT 210.760 189.010 217.505 189.150 ;
        RECT 191.455 188.625 191.745 188.855 ;
        RECT 194.200 188.810 194.520 188.870 ;
        RECT 197.055 188.810 197.195 188.965 ;
        RECT 210.760 188.950 211.080 189.010 ;
        RECT 217.215 188.965 217.505 189.010 ;
        RECT 225.020 189.150 225.340 189.210 ;
        RECT 227.335 189.150 227.625 189.195 ;
        RECT 225.020 189.010 227.625 189.150 ;
        RECT 225.020 188.950 225.340 189.010 ;
        RECT 227.335 188.965 227.625 189.010 ;
        RECT 228.240 188.950 228.560 189.210 ;
        RECT 229.160 189.150 229.480 189.210 ;
        RECT 230.095 189.150 230.385 189.195 ;
        RECT 232.395 189.150 232.685 189.195 ;
        RECT 229.160 189.010 230.385 189.150 ;
        RECT 229.160 188.950 229.480 189.010 ;
        RECT 230.095 188.965 230.385 189.010 ;
        RECT 230.630 189.010 232.685 189.150 ;
        RECT 194.200 188.670 197.195 188.810 ;
        RECT 229.620 188.810 229.940 188.870 ;
        RECT 230.630 188.810 230.770 189.010 ;
        RECT 232.395 188.965 232.685 189.010 ;
        RECT 233.775 188.965 234.065 189.195 ;
        RECT 229.620 188.670 230.770 188.810 ;
        RECT 231.000 188.810 231.320 188.870 ;
        RECT 233.850 188.810 233.990 188.965 ;
        RECT 231.000 188.670 233.990 188.810 ;
        RECT 187.300 188.470 187.620 188.530 ;
        RECT 186.010 188.330 187.620 188.470 ;
        RECT 187.300 188.270 187.620 188.330 ;
        RECT 188.235 188.470 188.525 188.515 ;
        RECT 191.530 188.470 191.670 188.625 ;
        RECT 194.200 188.610 194.520 188.670 ;
        RECT 229.620 188.610 229.940 188.670 ;
        RECT 231.000 188.610 231.320 188.670 ;
        RECT 188.235 188.330 191.670 188.470 ;
        RECT 198.355 188.470 198.645 188.515 ;
        RECT 199.720 188.470 200.040 188.530 ;
        RECT 198.355 188.330 200.040 188.470 ;
        RECT 188.235 188.285 188.525 188.330 ;
        RECT 198.355 188.285 198.645 188.330 ;
        RECT 199.720 188.270 200.040 188.330 ;
        RECT 227.320 188.470 227.640 188.530 ;
        RECT 231.475 188.470 231.765 188.515 ;
        RECT 227.320 188.330 231.765 188.470 ;
        RECT 227.320 188.270 227.640 188.330 ;
        RECT 231.475 188.285 231.765 188.330 ;
        RECT 149.905 185.540 150.865 185.770 ;
        RECT 151.195 185.540 152.155 185.770 ;
        RECT 152.845 185.165 155.165 187.965 ;
        RECT 165.150 187.650 239.210 188.130 ;
        RECT 167.980 187.250 168.300 187.510 ;
        RECT 168.440 187.450 168.760 187.510 ;
        RECT 172.135 187.450 172.425 187.495 ;
        RECT 168.440 187.310 172.425 187.450 ;
        RECT 168.440 187.250 168.760 187.310 ;
        RECT 172.135 187.265 172.425 187.310 ;
        RECT 175.815 187.450 176.105 187.495 ;
        RECT 176.260 187.450 176.580 187.510 ;
        RECT 180.860 187.450 181.180 187.510 ;
        RECT 175.815 187.310 181.180 187.450 ;
        RECT 175.815 187.265 176.105 187.310 ;
        RECT 176.260 187.250 176.580 187.310 ;
        RECT 180.860 187.250 181.180 187.310 ;
        RECT 182.240 187.250 182.560 187.510 ;
        RECT 183.635 187.450 183.925 187.495 ;
        RECT 186.380 187.450 186.700 187.510 ;
        RECT 183.635 187.310 186.700 187.450 ;
        RECT 183.635 187.265 183.925 187.310 ;
        RECT 186.380 187.250 186.700 187.310 ;
        RECT 189.140 187.450 189.460 187.510 ;
        RECT 193.740 187.450 194.060 187.510 ;
        RECT 189.140 187.310 194.060 187.450 ;
        RECT 189.140 187.250 189.460 187.310 ;
        RECT 193.740 187.250 194.060 187.310 ;
        RECT 201.115 187.265 201.405 187.495 ;
        RECT 208.015 187.450 208.305 187.495 ;
        RECT 208.920 187.450 209.240 187.510 ;
        RECT 208.015 187.310 209.240 187.450 ;
        RECT 208.015 187.265 208.305 187.310 ;
        RECT 179.940 187.110 180.260 187.170 ;
        RECT 168.530 186.970 180.260 187.110 ;
        RECT 168.530 186.815 168.670 186.970 ;
        RECT 179.940 186.910 180.260 186.970 ;
        RECT 180.400 186.910 180.720 187.170 ;
        RECT 184.540 187.110 184.860 187.170 ;
        RECT 186.840 187.110 187.160 187.170 ;
        RECT 184.540 186.970 187.160 187.110 ;
        RECT 184.540 186.910 184.860 186.970 ;
        RECT 186.840 186.910 187.160 186.970 ;
        RECT 189.600 187.110 189.920 187.170 ;
        RECT 189.600 186.970 198.575 187.110 ;
        RECT 189.600 186.910 189.920 186.970 ;
        RECT 167.075 186.585 167.365 186.815 ;
        RECT 168.455 186.585 168.745 186.815 ;
        RECT 168.900 186.770 169.220 186.830 ;
        RECT 169.835 186.770 170.125 186.815 ;
        RECT 168.900 186.630 170.125 186.770 ;
        RECT 167.150 185.750 167.290 186.585 ;
        RECT 168.900 186.570 169.220 186.630 ;
        RECT 169.835 186.585 170.125 186.630 ;
        RECT 170.280 186.770 170.600 186.830 ;
        RECT 173.515 186.770 173.805 186.815 ;
        RECT 170.280 186.630 173.805 186.770 ;
        RECT 170.280 186.570 170.600 186.630 ;
        RECT 173.515 186.585 173.805 186.630 ;
        RECT 175.800 186.770 176.120 186.830 ;
        RECT 176.275 186.770 176.565 186.815 ;
        RECT 175.800 186.630 176.565 186.770 ;
        RECT 175.800 186.570 176.120 186.630 ;
        RECT 176.275 186.585 176.565 186.630 ;
        RECT 177.195 186.770 177.485 186.815 ;
        RECT 177.640 186.770 177.960 186.830 ;
        RECT 177.195 186.630 177.960 186.770 ;
        RECT 177.195 186.585 177.485 186.630 ;
        RECT 177.640 186.570 177.960 186.630 ;
        RECT 178.115 186.585 178.405 186.815 ;
        RECT 179.495 186.770 179.785 186.815 ;
        RECT 180.860 186.770 181.180 186.830 ;
        RECT 179.495 186.630 181.180 186.770 ;
        RECT 179.495 186.585 179.785 186.630 ;
        RECT 167.520 186.430 167.840 186.490 ;
        RECT 178.190 186.430 178.330 186.585 ;
        RECT 180.860 186.570 181.180 186.630 ;
        RECT 181.335 186.770 181.625 186.815 ;
        RECT 182.240 186.770 182.560 186.830 ;
        RECT 181.335 186.630 182.560 186.770 ;
        RECT 181.335 186.585 181.625 186.630 ;
        RECT 182.240 186.570 182.560 186.630 ;
        RECT 182.715 186.770 183.005 186.815 ;
        RECT 183.620 186.770 183.940 186.830 ;
        RECT 182.715 186.630 183.940 186.770 ;
        RECT 182.715 186.585 183.005 186.630 ;
        RECT 183.620 186.570 183.940 186.630 ;
        RECT 185.000 186.570 185.320 186.830 ;
        RECT 185.475 186.770 185.765 186.815 ;
        RECT 185.920 186.770 186.240 186.830 ;
        RECT 185.475 186.630 186.240 186.770 ;
        RECT 185.475 186.585 185.765 186.630 ;
        RECT 185.920 186.570 186.240 186.630 ;
        RECT 187.760 186.570 188.080 186.830 ;
        RECT 189.140 186.570 189.460 186.830 ;
        RECT 190.060 186.770 190.380 186.830 ;
        RECT 190.535 186.770 190.825 186.815 ;
        RECT 190.060 186.630 190.825 186.770 ;
        RECT 190.060 186.570 190.380 186.630 ;
        RECT 190.535 186.585 190.825 186.630 ;
        RECT 191.440 186.770 191.760 186.830 ;
        RECT 191.915 186.770 192.205 186.815 ;
        RECT 191.440 186.630 192.205 186.770 ;
        RECT 191.440 186.570 191.760 186.630 ;
        RECT 191.915 186.585 192.205 186.630 ;
        RECT 193.740 186.570 194.060 186.830 ;
        RECT 194.295 186.815 194.435 186.970 ;
        RECT 198.435 186.830 198.575 186.970 ;
        RECT 199.720 186.910 200.040 187.170 ;
        RECT 201.190 187.110 201.330 187.265 ;
        RECT 208.920 187.250 209.240 187.310 ;
        RECT 209.380 187.450 209.700 187.510 ;
        RECT 225.020 187.450 225.340 187.510 ;
        RECT 209.380 187.310 225.340 187.450 ;
        RECT 209.380 187.250 209.700 187.310 ;
        RECT 225.020 187.250 225.340 187.310 ;
        RECT 231.935 187.450 232.225 187.495 ;
        RECT 232.380 187.450 232.700 187.510 ;
        RECT 231.935 187.310 232.700 187.450 ;
        RECT 231.935 187.265 232.225 187.310 ;
        RECT 232.380 187.250 232.700 187.310 ;
        RECT 234.695 187.450 234.985 187.495 ;
        RECT 236.060 187.450 236.380 187.510 ;
        RECT 234.695 187.310 236.380 187.450 ;
        RECT 234.695 187.265 234.985 187.310 ;
        RECT 236.060 187.250 236.380 187.310 ;
        RECT 210.760 187.110 211.080 187.170 ;
        RECT 201.190 186.970 211.080 187.110 ;
        RECT 210.760 186.910 211.080 186.970 ;
        RECT 211.220 187.110 211.540 187.170 ;
        RECT 218.120 187.110 218.440 187.170 ;
        RECT 219.960 187.110 220.280 187.170 ;
        RECT 224.120 187.110 224.410 187.155 ;
        RECT 229.640 187.110 229.930 187.155 ;
        RECT 230.560 187.110 230.850 187.155 ;
        RECT 211.220 186.970 213.750 187.110 ;
        RECT 211.220 186.910 211.540 186.970 ;
        RECT 194.220 186.585 194.510 186.815 ;
        RECT 195.120 186.570 195.440 186.830 ;
        RECT 196.040 186.815 196.360 186.830 ;
        RECT 195.595 186.585 195.885 186.815 ;
        RECT 196.040 186.585 196.370 186.815 ;
        RECT 197.895 186.770 198.185 186.815 ;
        RECT 196.590 186.630 198.185 186.770 ;
        RECT 167.520 186.290 178.330 186.430 ;
        RECT 192.360 186.430 192.680 186.490 ;
        RECT 195.670 186.430 195.810 186.585 ;
        RECT 196.040 186.570 196.360 186.585 ;
        RECT 192.360 186.290 195.810 186.430 ;
        RECT 167.520 186.230 167.840 186.290 ;
        RECT 192.360 186.230 192.680 186.290 ;
        RECT 169.375 186.090 169.665 186.135 ;
        RECT 178.100 186.090 178.420 186.150 ;
        RECT 186.855 186.090 187.145 186.135 ;
        RECT 169.375 185.950 178.420 186.090 ;
        RECT 169.375 185.905 169.665 185.950 ;
        RECT 178.100 185.890 178.420 185.950 ;
        RECT 178.650 185.950 187.145 186.090 ;
        RECT 169.820 185.750 170.140 185.810 ;
        RECT 167.150 185.610 170.140 185.750 ;
        RECT 169.820 185.550 170.140 185.610 ;
        RECT 170.740 185.550 171.060 185.810 ;
        RECT 176.720 185.750 177.040 185.810 ;
        RECT 178.650 185.750 178.790 185.950 ;
        RECT 186.855 185.905 187.145 185.950 ;
        RECT 193.740 186.090 194.060 186.150 ;
        RECT 196.590 186.090 196.730 186.630 ;
        RECT 197.895 186.585 198.185 186.630 ;
        RECT 198.340 186.570 198.660 186.830 ;
        RECT 199.260 186.570 199.580 186.830 ;
        RECT 200.180 186.815 200.500 186.830 ;
        RECT 200.180 186.770 200.510 186.815 ;
        RECT 200.180 186.630 200.695 186.770 ;
        RECT 200.180 186.585 200.510 186.630 ;
        RECT 200.180 186.570 200.500 186.585 ;
        RECT 202.480 186.570 202.800 186.830 ;
        RECT 208.935 186.585 209.225 186.815 ;
        RECT 196.960 186.430 197.280 186.490 ;
        RECT 209.010 186.430 209.150 186.585 ;
        RECT 210.300 186.570 210.620 186.830 ;
        RECT 211.695 186.585 211.985 186.815 ;
        RECT 196.960 186.290 209.150 186.430 ;
        RECT 196.960 186.230 197.280 186.290 ;
        RECT 209.840 186.230 210.160 186.490 ;
        RECT 193.740 185.950 196.730 186.090 ;
        RECT 198.800 186.090 199.120 186.150 ;
        RECT 201.575 186.090 201.865 186.135 ;
        RECT 198.800 185.950 201.865 186.090 ;
        RECT 193.740 185.890 194.060 185.950 ;
        RECT 198.800 185.890 199.120 185.950 ;
        RECT 201.575 185.905 201.865 185.950 ;
        RECT 207.080 186.090 207.400 186.150 ;
        RECT 210.775 186.090 211.065 186.135 ;
        RECT 211.770 186.090 211.910 186.585 ;
        RECT 213.060 186.570 213.380 186.830 ;
        RECT 213.610 186.815 213.750 186.970 ;
        RECT 218.120 186.970 219.270 187.110 ;
        RECT 218.120 186.910 218.440 186.970 ;
        RECT 213.535 186.585 213.825 186.815 ;
        RECT 214.915 186.585 215.205 186.815 ;
        RECT 215.360 186.770 215.680 186.830 ;
        RECT 217.215 186.770 217.505 186.815 ;
        RECT 215.360 186.630 217.505 186.770 ;
        RECT 212.140 186.230 212.460 186.490 ;
        RECT 212.600 186.430 212.920 186.490 ;
        RECT 214.990 186.430 215.130 186.585 ;
        RECT 215.360 186.570 215.680 186.630 ;
        RECT 217.215 186.585 217.505 186.630 ;
        RECT 218.580 186.570 218.900 186.830 ;
        RECT 219.130 186.770 219.270 186.970 ;
        RECT 219.960 186.970 221.570 187.110 ;
        RECT 219.960 186.910 220.280 186.970 ;
        RECT 221.430 186.815 221.570 186.970 ;
        RECT 224.120 186.970 230.850 187.110 ;
        RECT 224.120 186.925 224.410 186.970 ;
        RECT 229.640 186.925 229.930 186.970 ;
        RECT 230.560 186.925 230.850 186.970 ;
        RECT 227.780 186.815 228.100 186.830 ;
        RECT 220.895 186.770 221.185 186.815 ;
        RECT 219.130 186.630 221.185 186.770 ;
        RECT 220.895 186.585 221.185 186.630 ;
        RECT 221.355 186.585 221.645 186.815 ;
        RECT 225.040 186.770 225.330 186.815 ;
        RECT 226.880 186.770 227.170 186.815 ;
        RECT 225.040 186.630 227.170 186.770 ;
        RECT 225.040 186.585 225.330 186.630 ;
        RECT 226.880 186.585 227.170 186.630 ;
        RECT 227.780 186.585 228.210 186.815 ;
        RECT 229.225 186.770 229.515 186.815 ;
        RECT 231.065 186.770 231.355 186.815 ;
        RECT 229.225 186.630 231.355 186.770 ;
        RECT 229.225 186.585 229.515 186.630 ;
        RECT 231.065 186.585 231.355 186.630 ;
        RECT 232.395 186.770 232.685 186.815 ;
        RECT 232.840 186.770 233.160 186.830 ;
        RECT 232.395 186.630 233.160 186.770 ;
        RECT 232.395 186.585 232.685 186.630 ;
        RECT 227.780 186.570 228.100 186.585 ;
        RECT 232.840 186.570 233.160 186.630 ;
        RECT 233.760 186.570 234.080 186.830 ;
        RECT 236.060 186.570 236.380 186.830 ;
        RECT 222.735 186.430 223.025 186.475 ;
        RECT 212.600 186.290 215.130 186.430 ;
        RECT 218.210 186.290 223.025 186.430 ;
        RECT 212.600 186.230 212.920 186.290 ;
        RECT 207.080 185.950 211.065 186.090 ;
        RECT 207.080 185.890 207.400 185.950 ;
        RECT 210.775 185.905 211.065 185.950 ;
        RECT 211.310 185.950 211.910 186.090 ;
        RECT 212.230 186.090 212.370 186.230 ;
        RECT 218.210 186.135 218.350 186.290 ;
        RECT 222.735 186.245 223.025 186.290 ;
        RECT 223.655 186.245 223.945 186.475 ;
        RECT 212.230 185.950 217.890 186.090 ;
        RECT 176.720 185.610 178.790 185.750 ;
        RECT 176.720 185.550 177.040 185.610 ;
        RECT 184.080 185.550 184.400 185.810 ;
        RECT 186.380 185.550 186.700 185.810 ;
        RECT 187.300 185.750 187.620 185.810 ;
        RECT 188.235 185.750 188.525 185.795 ;
        RECT 187.300 185.610 188.525 185.750 ;
        RECT 187.300 185.550 187.620 185.610 ;
        RECT 188.235 185.565 188.525 185.610 ;
        RECT 188.680 185.750 189.000 185.810 ;
        RECT 189.615 185.750 189.905 185.795 ;
        RECT 188.680 185.610 189.905 185.750 ;
        RECT 188.680 185.550 189.000 185.610 ;
        RECT 189.615 185.565 189.905 185.610 ;
        RECT 192.820 185.550 193.140 185.810 ;
        RECT 196.975 185.750 197.265 185.795 ;
        RECT 209.380 185.750 209.700 185.810 ;
        RECT 196.975 185.610 209.700 185.750 ;
        RECT 196.975 185.565 197.265 185.610 ;
        RECT 209.380 185.550 209.700 185.610 ;
        RECT 209.840 185.750 210.160 185.810 ;
        RECT 211.310 185.750 211.450 185.950 ;
        RECT 209.840 185.610 211.450 185.750 ;
        RECT 211.680 185.750 212.000 185.810 ;
        RECT 212.155 185.750 212.445 185.795 ;
        RECT 211.680 185.610 212.445 185.750 ;
        RECT 209.840 185.550 210.160 185.610 ;
        RECT 211.680 185.550 212.000 185.610 ;
        RECT 212.155 185.565 212.445 185.610 ;
        RECT 214.455 185.750 214.745 185.795 ;
        RECT 214.900 185.750 215.220 185.810 ;
        RECT 214.455 185.610 215.220 185.750 ;
        RECT 214.455 185.565 214.745 185.610 ;
        RECT 214.900 185.550 215.220 185.610 ;
        RECT 215.835 185.750 216.125 185.795 ;
        RECT 217.200 185.750 217.520 185.810 ;
        RECT 215.835 185.610 217.520 185.750 ;
        RECT 217.750 185.750 217.890 185.950 ;
        RECT 218.135 185.905 218.425 186.135 ;
        RECT 219.975 186.090 220.265 186.135 ;
        RECT 218.670 185.950 220.265 186.090 ;
        RECT 218.670 185.750 218.810 185.950 ;
        RECT 219.975 185.905 220.265 185.950 ;
        RECT 220.420 186.090 220.740 186.150 ;
        RECT 223.730 186.090 223.870 186.245 ;
        RECT 227.320 186.230 227.640 186.490 ;
        RECT 228.715 186.430 229.005 186.475 ;
        RECT 228.715 186.290 230.770 186.430 ;
        RECT 228.715 186.245 229.005 186.290 ;
        RECT 220.420 185.950 223.870 186.090 ;
        RECT 225.480 186.090 225.800 186.150 ;
        RECT 225.955 186.090 226.245 186.135 ;
        RECT 225.480 185.950 226.245 186.090 ;
        RECT 220.420 185.890 220.740 185.950 ;
        RECT 225.480 185.890 225.800 185.950 ;
        RECT 225.955 185.905 226.245 185.950 ;
        RECT 226.915 186.090 227.205 186.135 ;
        RECT 230.145 186.090 230.435 186.135 ;
        RECT 226.915 185.950 230.435 186.090 ;
        RECT 230.630 186.090 230.770 186.290 ;
        RECT 231.920 186.090 232.240 186.150 ;
        RECT 230.630 185.950 232.240 186.090 ;
        RECT 226.915 185.905 227.205 185.950 ;
        RECT 230.145 185.905 230.435 185.950 ;
        RECT 231.920 185.890 232.240 185.950 ;
        RECT 217.750 185.610 218.810 185.750 ;
        RECT 215.835 185.565 216.125 185.610 ;
        RECT 217.200 185.550 217.520 185.610 ;
        RECT 219.500 185.550 219.820 185.810 ;
        RECT 222.260 185.550 222.580 185.810 ;
        RECT 229.160 185.750 229.480 185.810 ;
        RECT 232.855 185.750 233.145 185.795 ;
        RECT 229.160 185.610 233.145 185.750 ;
        RECT 229.160 185.550 229.480 185.610 ;
        RECT 232.855 185.565 233.145 185.610 ;
        RECT 235.140 185.550 235.460 185.810 ;
        RECT 108.515 184.765 155.165 185.165 ;
        RECT 165.150 184.930 239.210 185.410 ;
        RECT 167.520 184.530 167.840 184.790 ;
        RECT 168.455 184.730 168.745 184.775 ;
        RECT 168.900 184.730 169.220 184.790 ;
        RECT 168.455 184.590 169.220 184.730 ;
        RECT 168.455 184.545 168.745 184.590 ;
        RECT 168.900 184.530 169.220 184.590 ;
        RECT 169.835 184.730 170.125 184.775 ;
        RECT 172.120 184.730 172.440 184.790 ;
        RECT 169.835 184.590 172.440 184.730 ;
        RECT 169.835 184.545 170.125 184.590 ;
        RECT 172.120 184.530 172.440 184.590 ;
        RECT 177.655 184.730 177.945 184.775 ;
        RECT 178.560 184.730 178.880 184.790 ;
        RECT 177.655 184.590 178.880 184.730 ;
        RECT 177.655 184.545 177.945 184.590 ;
        RECT 178.560 184.530 178.880 184.590 ;
        RECT 185.015 184.730 185.305 184.775 ;
        RECT 186.840 184.730 187.160 184.790 ;
        RECT 185.015 184.590 187.160 184.730 ;
        RECT 185.015 184.545 185.305 184.590 ;
        RECT 186.840 184.530 187.160 184.590 ;
        RECT 187.315 184.730 187.605 184.775 ;
        RECT 192.375 184.730 192.665 184.775 ;
        RECT 193.280 184.730 193.600 184.790 ;
        RECT 187.315 184.590 191.235 184.730 ;
        RECT 187.315 184.545 187.605 184.590 ;
        RECT 176.260 184.390 176.580 184.450 ;
        RECT 181.795 184.390 182.085 184.435 ;
        RECT 191.095 184.390 191.235 184.590 ;
        RECT 192.375 184.590 193.600 184.730 ;
        RECT 192.375 184.545 192.665 184.590 ;
        RECT 193.280 184.530 193.600 184.590 ;
        RECT 197.420 184.730 197.740 184.790 ;
        RECT 202.480 184.730 202.800 184.790 ;
        RECT 211.220 184.730 211.540 184.790 ;
        RECT 197.420 184.590 202.800 184.730 ;
        RECT 197.420 184.530 197.740 184.590 ;
        RECT 202.480 184.530 202.800 184.590 ;
        RECT 210.620 184.590 211.540 184.730 ;
        RECT 191.900 184.390 192.220 184.450 ;
        RECT 200.195 184.390 200.485 184.435 ;
        RECT 201.100 184.390 201.420 184.450 ;
        RECT 210.620 184.390 210.760 184.590 ;
        RECT 211.220 184.530 211.540 184.590 ;
        RECT 213.060 184.730 213.380 184.790 ;
        RECT 216.740 184.730 217.060 184.790 ;
        RECT 217.215 184.730 217.505 184.775 ;
        RECT 213.060 184.590 216.510 184.730 ;
        RECT 213.060 184.530 213.380 184.590 ;
        RECT 172.670 184.250 175.390 184.390 ;
        RECT 166.600 183.510 166.920 183.770 ;
        RECT 168.440 183.710 168.760 183.770 ;
        RECT 169.375 183.710 169.665 183.755 ;
        RECT 168.440 183.570 169.665 183.710 ;
        RECT 168.440 183.510 168.760 183.570 ;
        RECT 169.375 183.525 169.665 183.570 ;
        RECT 169.820 183.710 170.140 183.770 ;
        RECT 172.670 183.755 172.810 184.250 ;
        RECT 175.250 184.050 175.390 184.250 ;
        RECT 176.260 184.250 181.090 184.390 ;
        RECT 176.260 184.190 176.580 184.250 ;
        RECT 176.350 184.050 176.490 184.190 ;
        RECT 175.250 183.910 176.490 184.050 ;
        RECT 178.100 184.050 178.420 184.110 ;
        RECT 178.100 183.910 179.710 184.050 ;
        RECT 175.250 183.770 175.390 183.910 ;
        RECT 178.100 183.850 178.420 183.910 ;
        RECT 170.525 183.710 170.815 183.755 ;
        RECT 169.820 183.570 170.815 183.710 ;
        RECT 169.450 183.030 169.590 183.525 ;
        RECT 169.820 183.510 170.140 183.570 ;
        RECT 170.525 183.525 170.815 183.570 ;
        RECT 172.590 183.525 172.880 183.755 ;
        RECT 173.055 183.710 173.345 183.755 ;
        RECT 174.420 183.710 174.740 183.770 ;
        RECT 175.250 183.755 175.660 183.770 ;
        RECT 173.055 183.570 174.740 183.710 ;
        RECT 173.055 183.525 173.345 183.570 ;
        RECT 174.420 183.510 174.740 183.570 ;
        RECT 175.175 183.525 175.660 183.755 ;
        RECT 175.340 183.510 175.660 183.525 ;
        RECT 176.260 183.510 176.580 183.770 ;
        RECT 177.180 183.755 177.500 183.770 ;
        RECT 176.965 183.525 177.500 183.755 ;
        RECT 177.180 183.510 177.500 183.525 ;
        RECT 177.640 183.710 177.960 183.770 ;
        RECT 179.570 183.755 179.710 183.910 ;
        RECT 180.950 183.770 181.090 184.250 ;
        RECT 181.795 184.250 190.750 184.390 ;
        RECT 191.095 184.250 191.670 184.390 ;
        RECT 181.795 184.205 182.085 184.250 ;
        RECT 181.410 183.910 187.075 184.050 ;
        RECT 178.575 183.710 178.865 183.755 ;
        RECT 177.640 183.570 178.865 183.710 ;
        RECT 177.640 183.510 177.960 183.570 ;
        RECT 178.575 183.525 178.865 183.570 ;
        RECT 179.495 183.525 179.785 183.755 ;
        RECT 180.860 183.510 181.180 183.770 ;
        RECT 171.200 183.170 171.520 183.430 ;
        RECT 171.660 183.170 171.980 183.430 ;
        RECT 175.815 183.370 176.105 183.415 ;
        RECT 178.100 183.370 178.420 183.430 ;
        RECT 181.410 183.370 181.550 183.910 ;
        RECT 186.935 183.770 187.075 183.910 ;
        RECT 182.240 183.710 182.560 183.770 ;
        RECT 182.715 183.710 183.005 183.755 ;
        RECT 182.240 183.570 183.005 183.710 ;
        RECT 182.240 183.510 182.560 183.570 ;
        RECT 182.715 183.525 183.005 183.570 ;
        RECT 184.080 183.510 184.400 183.770 ;
        RECT 184.540 183.510 184.860 183.770 ;
        RECT 186.380 183.755 186.700 183.770 ;
        RECT 186.340 183.710 186.700 183.755 ;
        RECT 186.185 183.570 186.700 183.710 ;
        RECT 186.340 183.525 186.700 183.570 ;
        RECT 186.380 183.510 186.700 183.525 ;
        RECT 186.845 183.755 187.165 183.770 ;
        RECT 189.600 183.760 189.920 183.770 ;
        RECT 189.510 183.755 189.920 183.760 ;
        RECT 186.845 183.525 187.375 183.755 ;
        RECT 188.695 183.525 188.985 183.755 ;
        RECT 189.435 183.525 189.920 183.755 ;
        RECT 190.610 183.710 190.750 184.250 ;
        RECT 191.530 184.050 191.670 184.250 ;
        RECT 191.900 184.250 198.570 184.390 ;
        RECT 191.900 184.190 192.220 184.250 ;
        RECT 192.360 184.050 192.680 184.110 ;
        RECT 191.530 183.910 192.680 184.050 ;
        RECT 192.360 183.850 192.680 183.910 ;
        RECT 194.200 184.050 194.520 184.110 ;
        RECT 195.135 184.050 195.425 184.095 ;
        RECT 194.200 183.910 195.425 184.050 ;
        RECT 194.200 183.850 194.520 183.910 ;
        RECT 195.135 183.865 195.425 183.910 ;
        RECT 191.020 183.710 191.310 183.755 ;
        RECT 190.610 183.570 191.310 183.710 ;
        RECT 191.020 183.525 191.310 183.570 ;
        RECT 193.740 183.710 194.060 183.770 ;
        RECT 197.880 183.755 198.200 183.770 ;
        RECT 196.975 183.710 197.265 183.755 ;
        RECT 193.740 183.570 197.265 183.710 ;
        RECT 186.845 183.510 187.165 183.525 ;
        RECT 175.815 183.230 178.420 183.370 ;
        RECT 175.815 183.185 176.105 183.230 ;
        RECT 178.100 183.170 178.420 183.230 ;
        RECT 180.090 183.230 181.550 183.370 ;
        RECT 181.780 183.370 182.100 183.430 ;
        RECT 184.630 183.370 184.770 183.510 ;
        RECT 181.780 183.230 184.770 183.370 ;
        RECT 185.460 183.370 185.780 183.430 ;
        RECT 188.770 183.370 188.910 183.525 ;
        RECT 189.600 183.510 189.920 183.525 ;
        RECT 193.740 183.510 194.060 183.570 ;
        RECT 196.975 183.525 197.265 183.570 ;
        RECT 197.715 183.525 198.200 183.755 ;
        RECT 198.430 183.710 198.570 184.250 ;
        RECT 200.195 184.250 201.420 184.390 ;
        RECT 200.195 184.205 200.485 184.250 ;
        RECT 201.100 184.190 201.420 184.250 ;
        RECT 208.090 184.250 210.760 184.390 ;
        RECT 212.195 184.390 212.485 184.435 ;
        RECT 215.425 184.390 215.715 184.435 ;
        RECT 212.195 184.250 215.715 184.390 ;
        RECT 216.370 184.390 216.510 184.590 ;
        RECT 216.740 184.590 217.505 184.730 ;
        RECT 216.740 184.530 217.060 184.590 ;
        RECT 217.215 184.545 217.505 184.590 ;
        RECT 220.050 184.590 228.930 184.730 ;
        RECT 219.040 184.390 219.360 184.450 ;
        RECT 216.370 184.250 219.360 184.390 ;
        RECT 208.090 184.095 208.230 184.250 ;
        RECT 212.195 184.205 212.485 184.250 ;
        RECT 215.425 184.205 215.715 184.250 ;
        RECT 219.040 184.190 219.360 184.250 ;
        RECT 208.015 183.865 208.305 184.095 ;
        RECT 209.380 184.050 209.700 184.110 ;
        RECT 211.235 184.050 211.525 184.095 ;
        RECT 209.380 183.910 211.525 184.050 ;
        RECT 209.380 183.850 209.700 183.910 ;
        RECT 211.235 183.865 211.525 183.910 ;
        RECT 211.680 184.050 212.000 184.110 ;
        RECT 213.060 184.095 213.380 184.110 ;
        RECT 212.615 184.050 212.905 184.095 ;
        RECT 211.680 183.910 212.905 184.050 ;
        RECT 211.680 183.850 212.000 183.910 ;
        RECT 212.615 183.865 212.905 183.910 ;
        RECT 213.060 183.865 213.490 184.095 ;
        RECT 213.060 183.850 213.380 183.865 ;
        RECT 213.980 183.850 214.300 184.110 ;
        RECT 214.900 184.050 215.220 184.110 ;
        RECT 215.820 184.050 216.140 184.110 ;
        RECT 220.050 184.095 220.190 184.590 ;
        RECT 221.340 184.390 221.660 184.450 ;
        RECT 223.195 184.390 223.485 184.435 ;
        RECT 221.340 184.250 223.485 184.390 ;
        RECT 221.340 184.190 221.660 184.250 ;
        RECT 223.195 184.205 223.485 184.250 ;
        RECT 224.155 184.390 224.445 184.435 ;
        RECT 227.385 184.390 227.675 184.435 ;
        RECT 224.155 184.250 227.675 184.390 ;
        RECT 228.790 184.390 228.930 184.590 ;
        RECT 229.160 184.530 229.480 184.790 ;
        RECT 230.080 184.730 230.400 184.790 ;
        RECT 230.080 184.590 232.150 184.730 ;
        RECT 230.080 184.530 230.400 184.590 ;
        RECT 230.540 184.390 230.860 184.450 ;
        RECT 228.790 184.250 230.860 184.390 ;
        RECT 224.155 184.205 224.445 184.250 ;
        RECT 227.385 184.205 227.675 184.250 ;
        RECT 230.540 184.190 230.860 184.250 ;
        RECT 231.475 184.205 231.765 184.435 ;
        RECT 232.010 184.390 232.150 184.590 ;
        RECT 234.220 184.530 234.540 184.790 ;
        RECT 232.010 184.250 235.370 184.390 ;
        RECT 214.900 183.910 216.140 184.050 ;
        RECT 214.900 183.850 215.220 183.910 ;
        RECT 215.820 183.850 216.140 183.910 ;
        RECT 219.975 183.865 220.265 184.095 ;
        RECT 224.560 183.850 224.880 184.110 ;
        RECT 225.265 184.050 225.555 184.095 ;
        RECT 231.550 184.050 231.690 184.205 ;
        RECT 225.265 183.910 231.690 184.050 ;
        RECT 225.265 183.865 225.555 183.910 ;
        RECT 199.300 183.710 199.590 183.755 ;
        RECT 198.430 183.570 199.590 183.710 ;
        RECT 199.300 183.525 199.590 183.570 ;
        RECT 200.640 183.710 200.960 183.770 ;
        RECT 202.035 183.710 202.325 183.755 ;
        RECT 200.640 183.570 202.325 183.710 ;
        RECT 197.880 183.510 198.200 183.525 ;
        RECT 200.640 183.510 200.960 183.570 ;
        RECT 202.035 183.525 202.325 183.570 ;
        RECT 203.415 183.525 203.705 183.755 ;
        RECT 206.635 183.710 206.925 183.755 ;
        RECT 208.460 183.710 208.780 183.770 ;
        RECT 206.635 183.570 208.780 183.710 ;
        RECT 206.635 183.525 206.925 183.570 ;
        RECT 185.460 183.230 188.910 183.370 ;
        RECT 180.090 183.030 180.230 183.230 ;
        RECT 181.780 183.170 182.100 183.230 ;
        RECT 185.460 183.170 185.780 183.230 ;
        RECT 190.060 183.170 190.380 183.430 ;
        RECT 190.535 183.370 190.825 183.415 ;
        RECT 196.500 183.370 196.820 183.430 ;
        RECT 190.535 183.230 191.210 183.370 ;
        RECT 190.535 183.185 190.825 183.230 ;
        RECT 191.070 183.090 191.210 183.230 ;
        RECT 193.370 183.230 196.820 183.370 ;
        RECT 169.450 182.890 180.230 183.030 ;
        RECT 180.400 183.030 180.720 183.090 ;
        RECT 183.635 183.030 183.925 183.075 ;
        RECT 180.400 182.890 183.925 183.030 ;
        RECT 180.400 182.830 180.720 182.890 ;
        RECT 183.635 182.845 183.925 182.890 ;
        RECT 190.980 182.830 191.300 183.090 ;
        RECT 191.915 183.030 192.205 183.075 ;
        RECT 193.370 183.030 193.510 183.230 ;
        RECT 196.500 183.170 196.820 183.230 ;
        RECT 198.340 183.170 198.660 183.430 ;
        RECT 198.815 183.185 199.105 183.415 ;
        RECT 203.490 183.370 203.630 183.525 ;
        RECT 208.460 183.510 208.780 183.570 ;
        RECT 208.935 183.525 209.225 183.755 ;
        RECT 210.320 183.710 210.610 183.755 ;
        RECT 212.160 183.710 212.450 183.755 ;
        RECT 210.320 183.570 212.450 183.710 ;
        RECT 210.320 183.525 210.610 183.570 ;
        RECT 212.160 183.525 212.450 183.570 ;
        RECT 214.505 183.710 214.795 183.755 ;
        RECT 216.345 183.710 216.635 183.755 ;
        RECT 214.505 183.570 216.635 183.710 ;
        RECT 214.505 183.525 214.795 183.570 ;
        RECT 216.345 183.525 216.635 183.570 ;
        RECT 209.010 183.370 209.150 183.525 ;
        RECT 217.660 183.510 217.980 183.770 ;
        RECT 220.895 183.525 221.185 183.755 ;
        RECT 222.280 183.710 222.570 183.755 ;
        RECT 224.120 183.710 224.410 183.755 ;
        RECT 222.280 183.570 224.410 183.710 ;
        RECT 222.280 183.525 222.570 183.570 ;
        RECT 224.120 183.525 224.410 183.570 ;
        RECT 199.810 183.230 203.630 183.370 ;
        RECT 203.950 183.230 209.150 183.370 ;
        RECT 209.400 183.370 209.690 183.415 ;
        RECT 214.920 183.370 215.210 183.415 ;
        RECT 215.840 183.370 216.130 183.415 ;
        RECT 220.970 183.370 221.110 183.525 ;
        RECT 225.940 183.510 226.260 183.770 ;
        RECT 226.465 183.710 226.755 183.755 ;
        RECT 228.305 183.710 228.595 183.755 ;
        RECT 226.465 183.570 228.595 183.710 ;
        RECT 226.465 183.525 226.755 183.570 ;
        RECT 228.305 183.525 228.595 183.570 ;
        RECT 229.160 183.710 229.480 183.770 ;
        RECT 231.015 183.710 231.305 183.755 ;
        RECT 229.160 183.570 231.305 183.710 ;
        RECT 229.160 183.510 229.480 183.570 ;
        RECT 231.015 183.525 231.305 183.570 ;
        RECT 232.395 183.525 232.685 183.755 ;
        RECT 233.775 183.710 234.065 183.755 ;
        RECT 234.220 183.710 234.540 183.770 ;
        RECT 235.230 183.755 235.370 184.250 ;
        RECT 233.775 183.570 234.540 183.710 ;
        RECT 233.775 183.525 234.065 183.570 ;
        RECT 209.400 183.230 216.130 183.370 ;
        RECT 191.915 182.890 193.510 183.030 ;
        RECT 193.740 183.030 194.060 183.090 ;
        RECT 194.215 183.030 194.505 183.075 ;
        RECT 193.740 182.890 194.505 183.030 ;
        RECT 191.915 182.845 192.205 182.890 ;
        RECT 193.740 182.830 194.060 182.890 ;
        RECT 194.215 182.845 194.505 182.890 ;
        RECT 194.660 182.830 194.980 183.090 ;
        RECT 195.580 183.030 195.900 183.090 ;
        RECT 198.890 183.030 199.030 183.185 ;
        RECT 199.810 183.090 199.950 183.230 ;
        RECT 195.580 182.890 199.030 183.030 ;
        RECT 195.580 182.830 195.900 182.890 ;
        RECT 199.720 182.830 200.040 183.090 ;
        RECT 201.100 182.830 201.420 183.090 ;
        RECT 201.560 183.030 201.880 183.090 ;
        RECT 202.495 183.030 202.785 183.075 ;
        RECT 201.560 182.890 202.785 183.030 ;
        RECT 201.560 182.830 201.880 182.890 ;
        RECT 202.495 182.845 202.785 182.890 ;
        RECT 203.400 183.030 203.720 183.090 ;
        RECT 203.950 183.030 204.090 183.230 ;
        RECT 209.400 183.185 209.690 183.230 ;
        RECT 214.920 183.185 215.210 183.230 ;
        RECT 215.840 183.185 216.130 183.230 ;
        RECT 218.210 183.230 221.110 183.370 ;
        RECT 221.360 183.370 221.650 183.415 ;
        RECT 226.880 183.370 227.170 183.415 ;
        RECT 227.800 183.370 228.090 183.415 ;
        RECT 232.470 183.370 232.610 183.525 ;
        RECT 234.220 183.510 234.540 183.570 ;
        RECT 235.155 183.525 235.445 183.755 ;
        RECT 236.535 183.525 236.825 183.755 ;
        RECT 221.360 183.230 228.090 183.370 ;
        RECT 203.400 182.890 204.090 183.030 ;
        RECT 207.555 183.030 207.845 183.075 ;
        RECT 218.210 183.030 218.350 183.230 ;
        RECT 221.360 183.185 221.650 183.230 ;
        RECT 226.880 183.185 227.170 183.230 ;
        RECT 227.800 183.185 228.090 183.230 ;
        RECT 228.330 183.230 232.610 183.370 ;
        RECT 233.300 183.370 233.620 183.430 ;
        RECT 236.610 183.370 236.750 183.525 ;
        RECT 233.300 183.230 236.750 183.370 ;
        RECT 207.555 182.890 218.350 183.030 ;
        RECT 218.595 183.030 218.885 183.075 ;
        RECT 224.100 183.030 224.420 183.090 ;
        RECT 218.595 182.890 224.420 183.030 ;
        RECT 203.400 182.830 203.720 182.890 ;
        RECT 207.555 182.845 207.845 182.890 ;
        RECT 218.595 182.845 218.885 182.890 ;
        RECT 224.100 182.830 224.420 182.890 ;
        RECT 224.560 183.030 224.880 183.090 ;
        RECT 228.330 183.030 228.470 183.230 ;
        RECT 233.300 183.170 233.620 183.230 ;
        RECT 224.560 182.890 228.470 183.030 ;
        RECT 224.560 182.830 224.880 182.890 ;
        RECT 230.080 182.830 230.400 183.090 ;
        RECT 232.840 182.830 233.160 183.090 ;
        RECT 235.600 182.830 235.920 183.090 ;
        RECT 63.895 181.400 64.595 182.400 ;
        RECT 77.595 182.370 78.595 182.605 ;
        RECT 77.595 181.195 78.595 181.430 ;
        RECT 80.185 181.400 81.755 182.400 ;
        RECT 83.345 182.370 84.345 182.605 ;
        RECT 83.345 181.195 84.345 181.430 ;
        RECT 97.345 181.400 98.045 182.400 ;
        RECT 64.175 180.965 80.135 181.195 ;
        RECT 81.805 180.965 97.765 181.195 ;
        RECT 77.595 180.730 78.595 180.965 ;
        RECT 83.345 180.730 84.345 180.965 ;
        RECT 98.485 180.110 155.900 182.710 ;
        RECT 165.150 182.210 239.210 182.690 ;
        RECT 168.455 182.010 168.745 182.055 ;
        RECT 169.820 182.010 170.140 182.070 ;
        RECT 168.455 181.870 170.140 182.010 ;
        RECT 168.455 181.825 168.745 181.870 ;
        RECT 169.820 181.810 170.140 181.870 ;
        RECT 171.660 182.010 171.980 182.070 ;
        RECT 172.135 182.010 172.425 182.055 ;
        RECT 171.660 181.870 172.425 182.010 ;
        RECT 171.660 181.810 171.980 181.870 ;
        RECT 172.135 181.825 172.425 181.870 ;
        RECT 173.040 181.810 173.360 182.070 ;
        RECT 173.975 182.010 174.265 182.055 ;
        RECT 175.800 182.010 176.120 182.070 ;
        RECT 173.975 181.870 176.120 182.010 ;
        RECT 173.975 181.825 174.265 181.870 ;
        RECT 175.800 181.810 176.120 181.870 ;
        RECT 176.720 182.010 177.040 182.070 ;
        RECT 179.940 182.010 180.260 182.070 ;
        RECT 176.720 181.870 180.260 182.010 ;
        RECT 176.720 181.810 177.040 181.870 ;
        RECT 179.940 181.810 180.260 181.870 ;
        RECT 186.380 181.810 186.700 182.070 ;
        RECT 186.855 182.010 187.145 182.055 ;
        RECT 188.220 182.010 188.540 182.070 ;
        RECT 186.855 181.870 188.540 182.010 ;
        RECT 186.855 181.825 187.145 181.870 ;
        RECT 188.220 181.810 188.540 181.870 ;
        RECT 188.680 181.810 189.000 182.070 ;
        RECT 192.360 182.010 192.680 182.070 ;
        RECT 194.675 182.010 194.965 182.055 ;
        RECT 195.120 182.010 195.440 182.070 ;
        RECT 192.360 181.870 193.360 182.010 ;
        RECT 192.360 181.810 192.680 181.870 ;
        RECT 173.130 181.670 173.270 181.810 ;
        RECT 171.750 181.530 173.270 181.670 ;
        RECT 174.435 181.670 174.725 181.715 ;
        RECT 178.560 181.670 178.880 181.730 ;
        RECT 174.435 181.530 178.880 181.670 ;
        RECT 167.060 181.130 167.380 181.390 ;
        RECT 169.375 181.330 169.665 181.375 ;
        RECT 169.375 181.190 170.510 181.330 ;
        RECT 169.375 181.145 169.665 181.190 ;
        RECT 167.995 180.650 168.285 180.695 ;
        RECT 169.360 180.650 169.680 180.710 ;
        RECT 167.995 180.510 169.680 180.650 ;
        RECT 170.370 180.650 170.510 181.190 ;
        RECT 170.740 181.130 171.060 181.390 ;
        RECT 171.750 181.375 171.890 181.530 ;
        RECT 174.435 181.485 174.725 181.530 ;
        RECT 178.560 181.470 178.880 181.530 ;
        RECT 181.320 181.670 181.640 181.730 ;
        RECT 189.155 181.670 189.445 181.715 ;
        RECT 181.320 181.530 184.310 181.670 ;
        RECT 181.320 181.470 181.640 181.530 ;
        RECT 171.735 181.145 172.025 181.375 ;
        RECT 176.735 181.330 177.025 181.375 ;
        RECT 177.180 181.330 177.500 181.390 ;
        RECT 176.735 181.190 177.500 181.330 ;
        RECT 176.735 181.145 177.025 181.190 ;
        RECT 177.180 181.130 177.500 181.190 ;
        RECT 178.115 181.145 178.405 181.375 ;
        RECT 170.830 180.990 170.970 181.130 ;
        RECT 175.355 180.990 175.645 181.035 ;
        RECT 177.640 180.990 177.960 181.050 ;
        RECT 170.830 180.850 177.960 180.990 ;
        RECT 178.190 180.990 178.330 181.145 ;
        RECT 179.020 181.130 179.340 181.390 ;
        RECT 180.415 181.330 180.705 181.375 ;
        RECT 180.860 181.330 181.180 181.390 ;
        RECT 180.415 181.190 181.180 181.330 ;
        RECT 180.415 181.145 180.705 181.190 ;
        RECT 180.860 181.130 181.180 181.190 ;
        RECT 181.780 181.130 182.100 181.390 ;
        RECT 182.715 181.330 183.005 181.375 ;
        RECT 183.160 181.330 183.480 181.390 ;
        RECT 184.170 181.375 184.310 181.530 ;
        RECT 189.155 181.530 190.750 181.670 ;
        RECT 189.155 181.485 189.445 181.530 ;
        RECT 190.610 181.390 190.750 181.530 ;
        RECT 182.715 181.190 183.480 181.330 ;
        RECT 182.715 181.145 183.005 181.190 ;
        RECT 183.160 181.130 183.480 181.190 ;
        RECT 184.095 181.145 184.385 181.375 ;
        RECT 185.460 181.130 185.780 181.390 ;
        RECT 188.220 181.330 188.540 181.390 ;
        RECT 186.930 181.250 189.830 181.330 ;
        RECT 186.700 181.190 189.830 181.250 ;
        RECT 181.870 180.990 182.010 181.130 ;
        RECT 186.700 181.110 187.070 181.190 ;
        RECT 188.220 181.130 188.540 181.190 ;
        RECT 186.700 180.990 186.840 181.110 ;
        RECT 189.690 181.035 189.830 181.190 ;
        RECT 190.520 181.130 190.840 181.390 ;
        RECT 190.980 181.330 191.300 181.390 ;
        RECT 193.220 181.375 193.360 181.870 ;
        RECT 194.675 181.870 195.440 182.010 ;
        RECT 194.675 181.825 194.965 181.870 ;
        RECT 195.120 181.810 195.440 181.870 ;
        RECT 198.340 182.010 198.660 182.070 ;
        RECT 198.815 182.010 199.105 182.055 ;
        RECT 198.340 181.870 199.105 182.010 ;
        RECT 198.340 181.810 198.660 181.870 ;
        RECT 198.815 181.825 199.105 181.870 ;
        RECT 200.180 182.010 200.500 182.070 ;
        RECT 200.655 182.010 200.945 182.055 ;
        RECT 200.180 181.870 200.945 182.010 ;
        RECT 200.180 181.810 200.500 181.870 ;
        RECT 200.655 181.825 200.945 181.870 ;
        RECT 205.255 182.010 205.545 182.055 ;
        RECT 210.300 182.010 210.620 182.070 ;
        RECT 205.255 181.870 210.620 182.010 ;
        RECT 205.255 181.825 205.545 181.870 ;
        RECT 210.300 181.810 210.620 181.870 ;
        RECT 222.720 182.010 223.040 182.070 ;
        RECT 229.160 182.010 229.480 182.070 ;
        RECT 222.720 181.870 229.480 182.010 ;
        RECT 222.720 181.810 223.040 181.870 ;
        RECT 229.160 181.810 229.480 181.870 ;
        RECT 232.380 182.010 232.700 182.070 ;
        RECT 236.535 182.010 236.825 182.055 ;
        RECT 232.380 181.870 236.825 182.010 ;
        RECT 232.380 181.810 232.700 181.870 ;
        RECT 236.535 181.825 236.825 181.870 ;
        RECT 196.975 181.670 197.265 181.715 ;
        RECT 201.100 181.670 201.420 181.730 ;
        RECT 206.160 181.670 206.480 181.730 ;
        RECT 196.975 181.530 201.420 181.670 ;
        RECT 196.975 181.485 197.265 181.530 ;
        RECT 201.100 181.470 201.420 181.530 ;
        RECT 204.410 181.530 206.480 181.670 ;
        RECT 192.375 181.330 192.665 181.375 ;
        RECT 190.980 181.190 192.665 181.330 ;
        RECT 190.980 181.130 191.300 181.190 ;
        RECT 192.375 181.145 192.665 181.190 ;
        RECT 193.145 181.330 193.435 181.375 ;
        RECT 193.145 181.190 194.890 181.330 ;
        RECT 193.145 181.145 193.435 181.190 ;
        RECT 178.190 180.850 186.840 180.990 ;
        RECT 189.615 180.990 189.905 181.035 ;
        RECT 194.200 180.990 194.520 181.050 ;
        RECT 189.615 180.850 194.520 180.990 ;
        RECT 194.750 180.990 194.890 181.190 ;
        RECT 196.500 181.130 196.820 181.390 ;
        RECT 202.480 181.330 202.800 181.390 ;
        RECT 204.410 181.375 204.550 181.530 ;
        RECT 206.160 181.470 206.480 181.530 ;
        RECT 208.480 181.670 208.770 181.715 ;
        RECT 214.000 181.670 214.290 181.715 ;
        RECT 214.920 181.670 215.210 181.715 ;
        RECT 208.480 181.530 215.210 181.670 ;
        RECT 208.480 181.485 208.770 181.530 ;
        RECT 214.000 181.485 214.290 181.530 ;
        RECT 214.920 181.485 215.210 181.530 ;
        RECT 218.600 181.670 218.890 181.715 ;
        RECT 224.120 181.670 224.410 181.715 ;
        RECT 225.040 181.670 225.330 181.715 ;
        RECT 218.600 181.530 225.330 181.670 ;
        RECT 218.600 181.485 218.890 181.530 ;
        RECT 224.120 181.485 224.410 181.530 ;
        RECT 225.040 181.485 225.330 181.530 ;
        RECT 228.260 181.670 228.550 181.715 ;
        RECT 233.780 181.670 234.070 181.715 ;
        RECT 234.700 181.670 234.990 181.715 ;
        RECT 228.260 181.530 234.990 181.670 ;
        RECT 228.260 181.485 228.550 181.530 ;
        RECT 233.780 181.485 234.070 181.530 ;
        RECT 234.700 181.485 234.990 181.530 ;
        RECT 202.955 181.330 203.245 181.375 ;
        RECT 202.480 181.190 203.245 181.330 ;
        RECT 202.480 181.130 202.800 181.190 ;
        RECT 202.955 181.145 203.245 181.190 ;
        RECT 204.335 181.145 204.625 181.375 ;
        RECT 205.240 181.330 205.560 181.390 ;
        RECT 205.715 181.330 206.005 181.375 ;
        RECT 209.400 181.330 209.690 181.375 ;
        RECT 211.240 181.330 211.530 181.375 ;
        RECT 205.240 181.190 206.005 181.330 ;
        RECT 205.240 181.130 205.560 181.190 ;
        RECT 205.715 181.145 206.005 181.190 ;
        RECT 206.710 181.190 208.690 181.330 ;
        RECT 197.435 180.990 197.725 181.035 ;
        RECT 194.750 180.850 197.725 180.990 ;
        RECT 175.355 180.805 175.645 180.850 ;
        RECT 177.640 180.790 177.960 180.850 ;
        RECT 179.110 180.710 179.250 180.850 ;
        RECT 189.615 180.805 189.905 180.850 ;
        RECT 194.200 180.790 194.520 180.850 ;
        RECT 197.435 180.805 197.725 180.850 ;
        RECT 197.880 180.990 198.200 181.050 ;
        RECT 201.115 180.990 201.405 181.035 ;
        RECT 197.880 180.850 201.405 180.990 ;
        RECT 170.370 180.510 174.650 180.650 ;
        RECT 167.995 180.465 168.285 180.510 ;
        RECT 169.360 180.450 169.680 180.510 ;
        RECT 174.510 180.370 174.650 180.510 ;
        RECT 179.020 180.450 179.340 180.710 ;
        RECT 180.400 180.650 180.720 180.710 ;
        RECT 190.980 180.650 191.300 180.710 ;
        RECT 180.400 180.510 191.300 180.650 ;
        RECT 197.510 180.650 197.650 180.805 ;
        RECT 197.880 180.790 198.200 180.850 ;
        RECT 201.115 180.805 201.405 180.850 ;
        RECT 202.020 180.790 202.340 181.050 ;
        RECT 206.710 180.990 206.850 181.190 ;
        RECT 202.570 180.850 206.850 180.990 ;
        RECT 202.570 180.650 202.710 180.850 ;
        RECT 207.080 180.790 207.400 181.050 ;
        RECT 208.015 180.805 208.305 181.035 ;
        RECT 208.550 180.990 208.690 181.190 ;
        RECT 209.400 181.190 211.530 181.330 ;
        RECT 209.400 181.145 209.690 181.190 ;
        RECT 211.240 181.145 211.530 181.190 ;
        RECT 213.585 181.330 213.875 181.375 ;
        RECT 215.425 181.330 215.715 181.375 ;
        RECT 213.585 181.190 215.715 181.330 ;
        RECT 213.585 181.145 213.875 181.190 ;
        RECT 215.425 181.145 215.715 181.190 ;
        RECT 217.200 181.130 217.520 181.390 ;
        RECT 222.260 181.375 222.580 181.390 ;
        RECT 219.520 181.330 219.810 181.375 ;
        RECT 221.360 181.330 221.650 181.375 ;
        RECT 219.520 181.190 221.650 181.330 ;
        RECT 219.520 181.145 219.810 181.190 ;
        RECT 221.360 181.145 221.650 181.190 ;
        RECT 222.260 181.145 222.690 181.375 ;
        RECT 223.705 181.330 223.995 181.375 ;
        RECT 225.545 181.330 225.835 181.375 ;
        RECT 223.705 181.190 225.835 181.330 ;
        RECT 223.705 181.145 223.995 181.190 ;
        RECT 225.545 181.145 225.835 181.190 ;
        RECT 229.180 181.330 229.470 181.375 ;
        RECT 231.020 181.330 231.310 181.375 ;
        RECT 231.565 181.330 231.855 181.375 ;
        RECT 229.180 181.190 231.310 181.330 ;
        RECT 231.550 181.310 231.855 181.330 ;
        RECT 229.180 181.145 229.470 181.190 ;
        RECT 231.020 181.145 231.310 181.190 ;
        RECT 231.460 181.145 231.855 181.310 ;
        RECT 222.260 181.130 222.580 181.145 ;
        RECT 231.460 181.050 231.780 181.145 ;
        RECT 232.840 181.130 233.160 181.390 ;
        RECT 233.365 181.330 233.655 181.375 ;
        RECT 235.205 181.330 235.495 181.375 ;
        RECT 237.455 181.330 237.745 181.375 ;
        RECT 233.365 181.190 235.495 181.330 ;
        RECT 233.365 181.145 233.655 181.190 ;
        RECT 235.205 181.145 235.495 181.190 ;
        RECT 235.690 181.190 237.745 181.330 ;
        RECT 210.315 180.990 210.605 181.035 ;
        RECT 208.550 180.850 210.605 180.990 ;
        RECT 197.510 180.510 202.710 180.650 ;
        RECT 203.875 180.650 204.165 180.695 ;
        RECT 208.090 180.650 208.230 180.805 ;
        RECT 209.470 180.710 209.610 180.850 ;
        RECT 210.315 180.805 210.605 180.850 ;
        RECT 211.680 180.790 212.000 181.050 ;
        RECT 212.140 181.035 212.460 181.050 ;
        RECT 212.140 180.805 212.570 181.035 ;
        RECT 212.140 180.790 212.460 180.805 ;
        RECT 213.060 180.790 213.380 181.050 ;
        RECT 218.135 180.990 218.425 181.035 ;
        RECT 214.990 180.850 218.425 180.990 ;
        RECT 203.875 180.510 208.230 180.650 ;
        RECT 180.400 180.450 180.720 180.510 ;
        RECT 190.980 180.450 191.300 180.510 ;
        RECT 203.875 180.465 204.165 180.510 ;
        RECT 209.380 180.450 209.700 180.710 ;
        RECT 211.275 180.650 211.565 180.695 ;
        RECT 214.505 180.650 214.795 180.695 ;
        RECT 211.275 180.510 214.795 180.650 ;
        RECT 211.275 180.465 211.565 180.510 ;
        RECT 214.505 180.465 214.795 180.510 ;
        RECT 174.420 180.310 174.740 180.370 ;
        RECT 175.340 180.310 175.660 180.370 ;
        RECT 174.420 180.170 175.660 180.310 ;
        RECT 174.420 180.110 174.740 180.170 ;
        RECT 175.340 180.110 175.660 180.170 ;
        RECT 177.640 180.110 177.960 180.370 ;
        RECT 181.335 180.310 181.625 180.355 ;
        RECT 184.540 180.310 184.860 180.370 ;
        RECT 181.335 180.170 184.860 180.310 ;
        RECT 181.335 180.125 181.625 180.170 ;
        RECT 184.540 180.110 184.860 180.170 ;
        RECT 185.015 180.310 185.305 180.355 ;
        RECT 191.900 180.310 192.220 180.370 ;
        RECT 185.015 180.170 192.220 180.310 ;
        RECT 185.015 180.125 185.305 180.170 ;
        RECT 191.900 180.110 192.220 180.170 ;
        RECT 193.295 180.310 193.585 180.355 ;
        RECT 195.580 180.310 195.900 180.370 ;
        RECT 193.295 180.170 195.900 180.310 ;
        RECT 193.295 180.125 193.585 180.170 ;
        RECT 195.580 180.110 195.900 180.170 ;
        RECT 206.635 180.310 206.925 180.355 ;
        RECT 214.990 180.310 215.130 180.850 ;
        RECT 218.135 180.805 218.425 180.850 ;
        RECT 221.800 180.790 222.120 181.050 ;
        RECT 223.180 180.790 223.500 181.050 ;
        RECT 224.100 180.990 224.420 181.050 ;
        RECT 226.875 180.990 227.165 181.035 ;
        RECT 224.100 180.850 227.165 180.990 ;
        RECT 224.100 180.790 224.420 180.850 ;
        RECT 226.875 180.805 227.165 180.850 ;
        RECT 227.780 180.790 228.100 181.050 ;
        RECT 232.380 181.035 232.700 181.050 ;
        RECT 232.165 180.805 232.700 181.035 ;
        RECT 232.380 180.790 232.700 180.805 ;
        RECT 216.280 180.450 216.600 180.710 ;
        RECT 217.200 180.650 217.520 180.710 ;
        RECT 220.435 180.650 220.725 180.695 ;
        RECT 217.200 180.510 220.725 180.650 ;
        RECT 217.200 180.450 217.520 180.510 ;
        RECT 220.435 180.465 220.725 180.510 ;
        RECT 221.395 180.650 221.685 180.695 ;
        RECT 224.625 180.650 224.915 180.695 ;
        RECT 225.480 180.650 225.800 180.710 ;
        RECT 230.095 180.650 230.385 180.695 ;
        RECT 221.395 180.510 224.915 180.650 ;
        RECT 221.395 180.465 221.685 180.510 ;
        RECT 224.625 180.465 224.915 180.510 ;
        RECT 225.110 180.510 230.385 180.650 ;
        RECT 206.635 180.170 215.130 180.310 ;
        RECT 220.510 180.310 220.650 180.465 ;
        RECT 225.110 180.310 225.250 180.510 ;
        RECT 225.480 180.450 225.800 180.510 ;
        RECT 230.095 180.465 230.385 180.510 ;
        RECT 231.055 180.650 231.345 180.695 ;
        RECT 234.285 180.650 234.575 180.695 ;
        RECT 231.055 180.510 234.575 180.650 ;
        RECT 231.055 180.465 231.345 180.510 ;
        RECT 234.285 180.465 234.575 180.510 ;
        RECT 220.510 180.170 225.250 180.310 ;
        RECT 206.635 180.125 206.925 180.170 ;
        RECT 226.400 180.110 226.720 180.370 ;
        RECT 227.780 180.310 228.100 180.370 ;
        RECT 235.690 180.310 235.830 181.190 ;
        RECT 237.455 181.145 237.745 181.190 ;
        RECT 236.075 180.990 236.365 181.035 ;
        RECT 236.520 180.990 236.840 181.050 ;
        RECT 236.075 180.850 236.840 180.990 ;
        RECT 236.075 180.805 236.365 180.850 ;
        RECT 236.520 180.790 236.840 180.850 ;
        RECT 227.780 180.170 235.830 180.310 ;
        RECT 227.780 180.110 228.100 180.170 ;
        RECT 77.595 179.815 78.595 180.050 ;
        RECT 83.345 179.815 84.345 180.050 ;
        RECT 64.175 179.585 80.135 179.815 ;
        RECT 81.805 179.585 97.765 179.815 ;
        RECT 63.895 178.380 64.595 179.380 ;
        RECT 77.595 179.350 78.595 179.585 ;
        RECT 77.595 178.175 78.595 178.410 ;
        RECT 80.185 178.380 81.755 179.380 ;
        RECT 83.345 179.350 84.345 179.585 ;
        RECT 83.345 178.175 84.345 178.410 ;
        RECT 97.345 178.380 98.045 179.380 ;
        RECT 64.175 177.945 80.135 178.175 ;
        RECT 81.805 177.945 97.765 178.175 ;
        RECT 77.595 177.710 78.595 177.945 ;
        RECT 83.345 177.710 84.345 177.945 ;
        RECT 77.595 176.795 78.595 177.030 ;
        RECT 83.345 176.795 84.345 177.030 ;
        RECT 64.175 176.565 80.135 176.795 ;
        RECT 81.805 176.565 97.765 176.795 ;
        RECT 63.895 175.360 64.595 176.360 ;
        RECT 77.595 176.330 78.595 176.565 ;
        RECT 77.595 175.155 78.595 175.390 ;
        RECT 80.185 175.360 81.755 176.360 ;
        RECT 83.345 176.330 84.345 176.565 ;
        RECT 83.345 175.155 84.345 175.390 ;
        RECT 97.345 175.360 98.045 176.360 ;
        RECT 64.175 174.925 80.135 175.155 ;
        RECT 81.805 174.925 97.765 175.155 ;
        RECT 77.595 174.690 78.595 174.925 ;
        RECT 83.345 174.690 84.345 174.925 ;
        RECT 64.175 173.545 80.135 173.775 ;
        RECT 81.805 173.545 97.765 173.775 ;
        RECT 63.895 172.340 64.125 173.340 ;
        RECT 80.185 172.340 81.755 173.340 ;
        RECT 97.815 172.340 98.045 173.340 ;
        RECT 64.175 171.905 80.135 172.135 ;
        RECT 81.805 171.905 97.765 172.135 ;
        RECT 98.485 171.445 100.480 180.110 ;
        RECT 62.865 160.555 100.480 171.445 ;
        RECT 5.910 143.155 58.705 143.745 ;
        RECT 5.910 140.725 23.785 143.155 ;
        RECT 24.505 143.045 25.505 143.155 ;
        RECT 24.255 142.435 57.645 142.665 ;
        RECT 24.255 141.275 24.485 142.435 ;
        RECT 28.015 141.965 29.015 142.435 ;
        RECT 32.545 141.275 32.775 142.435 ;
        RECT 36.305 141.965 37.305 142.435 ;
        RECT 40.835 141.275 41.065 142.435 ;
        RECT 44.595 141.965 45.595 142.435 ;
        RECT 49.125 141.275 49.355 142.435 ;
        RECT 52.885 141.965 53.885 142.435 ;
        RECT 57.415 141.275 57.645 142.435 ;
        RECT 24.535 140.885 32.495 141.115 ;
        RECT 32.825 140.885 40.785 141.115 ;
        RECT 41.115 140.885 49.075 141.115 ;
        RECT 49.405 140.885 57.365 141.115 ;
        RECT 5.910 139.725 24.955 140.725 ;
        RECT 32.545 139.725 32.775 140.725 ;
        RECT 40.835 139.725 41.065 140.725 ;
        RECT 49.125 139.725 49.355 140.725 ;
        RECT 56.545 139.725 57.645 140.725 ;
        RECT 5.910 139.175 23.785 139.725 ;
        RECT 24.535 139.335 32.495 139.565 ;
        RECT 32.825 139.335 40.785 139.565 ;
        RECT 41.115 139.335 49.075 139.565 ;
        RECT 49.405 139.335 57.365 139.565 ;
        RECT 5.910 138.175 24.955 139.175 ;
        RECT 32.545 138.175 32.775 139.175 ;
        RECT 40.835 138.175 41.065 139.175 ;
        RECT 49.125 138.175 49.355 139.175 ;
        RECT 53.035 138.175 57.645 139.175 ;
        RECT 5.910 137.925 23.785 138.175 ;
        RECT 5.910 137.075 9.990 137.925 ;
        RECT 11.145 137.465 11.845 137.535 ;
        RECT 14.080 137.465 14.780 137.535 ;
        RECT 15.370 137.465 16.070 137.535 ;
        RECT 18.305 137.465 19.005 137.535 ;
        RECT 11.015 137.235 11.975 137.465 ;
        RECT 13.950 137.235 14.910 137.465 ;
        RECT 15.240 137.235 16.200 137.465 ;
        RECT 18.175 137.235 19.135 137.465 ;
        RECT 5.910 136.075 10.965 137.075 ;
        RECT 12.025 136.925 12.255 137.075 ;
        RECT 11.990 136.225 12.290 136.925 ;
        RECT 12.025 136.075 12.255 136.225 ;
        RECT 5.910 135.225 9.990 136.075 ;
        RECT 13.670 135.825 13.900 137.075 ;
        RECT 14.960 136.925 15.190 137.075 ;
        RECT 16.250 136.925 16.480 137.075 ;
        RECT 14.925 136.225 15.225 136.925 ;
        RECT 16.215 136.225 16.515 136.925 ;
        RECT 14.960 136.075 15.190 136.225 ;
        RECT 16.250 136.075 16.480 136.225 ;
        RECT 13.435 135.525 14.135 135.825 ;
        RECT 17.895 135.225 18.125 137.075 ;
        RECT 19.185 136.775 19.415 137.075 ;
        RECT 19.150 136.075 19.450 136.775 ;
        RECT 20.160 135.745 23.785 137.925 ;
        RECT 24.535 137.785 32.495 138.015 ;
        RECT 32.825 137.785 40.785 138.015 ;
        RECT 41.115 137.785 49.075 138.015 ;
        RECT 49.405 137.785 57.365 138.015 ;
        RECT 24.255 136.465 24.485 137.625 ;
        RECT 28.015 136.465 29.015 136.935 ;
        RECT 32.545 136.465 32.775 137.625 ;
        RECT 36.305 136.465 37.305 136.935 ;
        RECT 40.835 136.465 41.065 137.625 ;
        RECT 44.595 136.465 45.595 136.935 ;
        RECT 49.125 136.465 49.355 137.625 ;
        RECT 52.885 136.465 53.885 136.935 ;
        RECT 57.415 136.465 57.645 137.625 ;
        RECT 24.255 136.235 57.645 136.465 ;
        RECT 24.505 135.745 25.505 135.855 ;
        RECT 58.115 135.745 58.705 143.155 ;
        RECT 20.160 135.225 58.705 135.745 ;
        RECT 5.910 132.225 58.705 135.225 ;
        RECT 62.865 139.455 69.970 160.555 ;
        RECT 71.220 157.040 89.820 159.315 ;
        RECT 71.220 142.990 73.495 157.040 ;
        RECT 76.385 157.030 77.215 157.040 ;
        RECT 80.105 157.030 80.935 157.040 ;
        RECT 83.825 157.030 84.655 157.040 ;
        RECT 74.940 154.420 86.100 155.595 ;
        RECT 74.940 153.050 76.115 154.420 ;
        RECT 76.385 153.310 77.215 154.140 ;
        RECT 77.485 153.050 79.835 154.420 ;
        RECT 80.105 153.310 80.935 154.140 ;
        RECT 81.205 153.050 83.555 154.420 ;
        RECT 83.825 153.310 84.655 154.140 ;
        RECT 84.925 153.050 86.100 154.420 ;
        RECT 74.940 150.700 86.100 153.050 ;
        RECT 74.940 149.330 76.115 150.700 ;
        RECT 76.385 149.590 77.215 150.420 ;
        RECT 77.485 149.330 79.835 150.700 ;
        RECT 80.105 149.590 80.935 150.420 ;
        RECT 81.205 149.330 83.555 150.700 ;
        RECT 83.825 149.590 84.655 150.420 ;
        RECT 84.925 149.330 86.100 150.700 ;
        RECT 74.940 146.980 86.100 149.330 ;
        RECT 74.940 145.610 76.115 146.980 ;
        RECT 76.385 145.870 77.215 146.700 ;
        RECT 77.485 145.610 79.835 146.980 ;
        RECT 80.105 145.870 80.935 146.700 ;
        RECT 81.205 145.610 83.555 146.980 ;
        RECT 83.825 145.870 84.655 146.700 ;
        RECT 84.925 145.610 86.100 146.980 ;
        RECT 74.940 144.435 86.100 145.610 ;
        RECT 87.545 142.990 89.820 157.040 ;
        RECT 71.220 140.715 89.820 142.990 ;
        RECT 91.070 139.455 100.480 160.555 ;
        RECT 101.935 176.325 152.755 178.210 ;
        RECT 101.935 174.870 114.420 176.325 ;
        RECT 115.200 175.635 118.030 176.165 ;
        RECT 119.820 175.635 122.650 176.165 ;
        RECT 124.440 175.635 127.270 176.165 ;
        RECT 129.060 175.635 131.890 176.165 ;
        RECT 133.680 175.635 136.510 176.165 ;
        RECT 138.300 175.635 141.130 176.165 ;
        RECT 142.920 175.635 145.750 176.165 ;
        RECT 147.540 175.635 150.370 176.165 ;
        RECT 114.920 174.870 115.150 175.475 ;
        RECT 101.935 172.215 115.185 174.870 ;
        RECT 101.935 162.685 103.025 172.215 ;
        RECT 103.715 171.610 104.675 171.840 ;
        RECT 105.005 171.610 105.965 171.840 ;
        RECT 103.435 170.840 103.665 171.450 ;
        RECT 103.400 168.540 103.700 170.840 ;
        RECT 103.435 163.450 103.665 168.540 ;
        RECT 104.725 167.140 104.955 171.450 ;
        RECT 106.015 170.840 106.245 171.450 ;
        RECT 105.980 168.540 106.280 170.840 ;
        RECT 104.690 164.840 104.990 167.140 ;
        RECT 104.725 163.450 104.955 164.840 ;
        RECT 106.015 163.450 106.245 168.540 ;
        RECT 103.715 163.060 104.675 163.290 ;
        RECT 105.005 163.060 105.965 163.290 ;
        RECT 103.715 162.990 104.415 163.060 ;
        RECT 105.265 162.990 105.965 163.060 ;
        RECT 106.655 162.685 107.055 172.215 ;
        RECT 110.685 172.070 115.185 172.215 ;
        RECT 107.745 171.610 108.705 171.840 ;
        RECT 109.035 171.610 109.995 171.840 ;
        RECT 107.465 170.840 107.695 171.450 ;
        RECT 107.430 168.540 107.730 170.840 ;
        RECT 107.465 163.450 107.695 168.540 ;
        RECT 108.755 167.140 108.985 171.450 ;
        RECT 110.045 170.840 110.275 171.450 ;
        RECT 110.010 168.540 110.310 170.840 ;
        RECT 108.720 164.840 109.020 167.140 ;
        RECT 108.755 163.450 108.985 164.840 ;
        RECT 110.045 163.450 110.275 168.540 ;
        RECT 110.685 166.625 114.420 172.070 ;
        RECT 114.920 167.475 115.150 172.070 ;
        RECT 115.710 170.895 115.940 175.475 ;
        RECT 116.500 174.870 116.730 175.475 ;
        RECT 116.465 172.070 116.765 174.870 ;
        RECT 115.675 168.095 115.975 170.895 ;
        RECT 115.710 167.475 115.940 168.095 ;
        RECT 116.500 167.475 116.730 172.070 ;
        RECT 117.290 170.895 117.520 175.475 ;
        RECT 118.080 174.870 118.310 175.475 ;
        RECT 119.540 174.870 119.770 175.475 ;
        RECT 118.045 172.070 118.345 174.870 ;
        RECT 119.505 172.070 119.805 174.870 ;
        RECT 117.255 168.095 117.555 170.895 ;
        RECT 117.290 167.475 117.520 168.095 ;
        RECT 118.080 167.475 118.310 172.070 ;
        RECT 119.540 167.475 119.770 172.070 ;
        RECT 120.330 170.895 120.560 175.475 ;
        RECT 121.120 174.870 121.350 175.475 ;
        RECT 121.085 172.070 121.385 174.870 ;
        RECT 120.295 168.095 120.595 170.895 ;
        RECT 120.330 167.475 120.560 168.095 ;
        RECT 121.120 167.475 121.350 172.070 ;
        RECT 121.910 170.895 122.140 175.475 ;
        RECT 122.700 174.870 122.930 175.475 ;
        RECT 124.160 174.870 124.390 175.475 ;
        RECT 122.665 172.070 122.965 174.870 ;
        RECT 124.125 172.070 124.425 174.870 ;
        RECT 121.875 168.095 122.175 170.895 ;
        RECT 121.910 167.475 122.140 168.095 ;
        RECT 122.700 167.475 122.930 172.070 ;
        RECT 124.160 167.475 124.390 172.070 ;
        RECT 124.950 170.895 125.180 175.475 ;
        RECT 125.740 174.870 125.970 175.475 ;
        RECT 125.705 172.070 126.005 174.870 ;
        RECT 124.915 168.095 125.215 170.895 ;
        RECT 124.950 167.475 125.180 168.095 ;
        RECT 125.740 167.475 125.970 172.070 ;
        RECT 126.530 170.895 126.760 175.475 ;
        RECT 127.320 174.870 127.550 175.475 ;
        RECT 128.780 174.870 129.010 175.475 ;
        RECT 127.285 172.070 127.585 174.870 ;
        RECT 128.745 172.070 129.045 174.870 ;
        RECT 126.495 168.095 126.795 170.895 ;
        RECT 126.530 167.475 126.760 168.095 ;
        RECT 127.320 167.475 127.550 172.070 ;
        RECT 128.780 167.475 129.010 172.070 ;
        RECT 129.570 170.895 129.800 175.475 ;
        RECT 130.360 174.870 130.590 175.475 ;
        RECT 130.325 172.070 130.625 174.870 ;
        RECT 129.535 168.095 129.835 170.895 ;
        RECT 129.570 167.475 129.800 168.095 ;
        RECT 130.360 167.475 130.590 172.070 ;
        RECT 131.150 170.895 131.380 175.475 ;
        RECT 131.940 174.870 132.170 175.475 ;
        RECT 133.400 174.870 133.630 175.475 ;
        RECT 131.905 172.070 132.205 174.870 ;
        RECT 133.365 172.070 133.665 174.870 ;
        RECT 131.115 168.095 131.415 170.895 ;
        RECT 131.150 167.475 131.380 168.095 ;
        RECT 131.940 167.475 132.170 172.070 ;
        RECT 133.400 167.475 133.630 172.070 ;
        RECT 134.190 170.895 134.420 175.475 ;
        RECT 134.980 174.870 135.210 175.475 ;
        RECT 134.945 172.070 135.245 174.870 ;
        RECT 134.155 168.095 134.455 170.895 ;
        RECT 134.190 167.475 134.420 168.095 ;
        RECT 134.980 167.475 135.210 172.070 ;
        RECT 135.770 170.895 136.000 175.475 ;
        RECT 136.560 174.870 136.790 175.475 ;
        RECT 138.020 174.870 138.250 175.475 ;
        RECT 136.525 172.070 136.825 174.870 ;
        RECT 137.985 172.070 138.285 174.870 ;
        RECT 135.735 168.095 136.035 170.895 ;
        RECT 135.770 167.475 136.000 168.095 ;
        RECT 136.560 167.475 136.790 172.070 ;
        RECT 138.020 167.475 138.250 172.070 ;
        RECT 138.810 170.895 139.040 175.475 ;
        RECT 139.600 174.870 139.830 175.475 ;
        RECT 139.565 172.070 139.865 174.870 ;
        RECT 138.775 168.095 139.075 170.895 ;
        RECT 138.810 167.475 139.040 168.095 ;
        RECT 139.600 167.475 139.830 172.070 ;
        RECT 140.390 170.895 140.620 175.475 ;
        RECT 141.180 174.870 141.410 175.475 ;
        RECT 142.640 174.870 142.870 175.475 ;
        RECT 141.145 172.070 141.445 174.870 ;
        RECT 142.605 172.070 142.905 174.870 ;
        RECT 140.355 168.095 140.655 170.895 ;
        RECT 140.390 167.475 140.620 168.095 ;
        RECT 141.180 167.475 141.410 172.070 ;
        RECT 142.640 167.475 142.870 172.070 ;
        RECT 143.430 170.895 143.660 175.475 ;
        RECT 144.220 174.870 144.450 175.475 ;
        RECT 144.185 172.070 144.485 174.870 ;
        RECT 143.395 168.095 143.695 170.895 ;
        RECT 143.430 167.475 143.660 168.095 ;
        RECT 144.220 167.475 144.450 172.070 ;
        RECT 145.010 170.895 145.240 175.475 ;
        RECT 145.800 174.870 146.030 175.475 ;
        RECT 147.260 174.870 147.490 175.475 ;
        RECT 145.765 172.070 146.065 174.870 ;
        RECT 147.225 172.070 147.525 174.870 ;
        RECT 144.975 168.095 145.275 170.895 ;
        RECT 145.010 167.475 145.240 168.095 ;
        RECT 145.800 167.475 146.030 172.070 ;
        RECT 147.260 167.475 147.490 172.070 ;
        RECT 148.050 170.895 148.280 175.475 ;
        RECT 148.840 174.870 149.070 175.475 ;
        RECT 148.805 172.070 149.105 174.870 ;
        RECT 148.015 168.095 148.315 170.895 ;
        RECT 148.050 167.475 148.280 168.095 ;
        RECT 148.840 167.475 149.070 172.070 ;
        RECT 149.630 170.895 149.860 175.475 ;
        RECT 150.420 174.870 150.650 175.475 ;
        RECT 150.385 172.070 150.685 174.870 ;
        RECT 149.595 168.095 149.895 170.895 ;
        RECT 149.630 167.475 149.860 168.095 ;
        RECT 150.420 167.475 150.650 172.070 ;
        RECT 115.200 167.085 115.660 167.315 ;
        RECT 115.990 167.085 116.450 167.315 ;
        RECT 116.780 167.085 117.240 167.315 ;
        RECT 117.570 167.085 118.030 167.315 ;
        RECT 119.820 167.085 120.280 167.315 ;
        RECT 120.610 167.085 121.070 167.315 ;
        RECT 121.400 167.085 121.860 167.315 ;
        RECT 122.190 167.085 122.650 167.315 ;
        RECT 124.440 167.085 124.900 167.315 ;
        RECT 125.230 167.085 125.690 167.315 ;
        RECT 126.020 167.085 126.480 167.315 ;
        RECT 126.810 167.085 127.270 167.315 ;
        RECT 129.060 167.085 129.520 167.315 ;
        RECT 129.850 167.085 130.310 167.315 ;
        RECT 130.640 167.085 131.100 167.315 ;
        RECT 131.430 167.085 131.890 167.315 ;
        RECT 133.680 167.085 134.140 167.315 ;
        RECT 134.470 167.085 134.930 167.315 ;
        RECT 135.260 167.085 135.720 167.315 ;
        RECT 136.050 167.085 136.510 167.315 ;
        RECT 138.300 167.085 138.760 167.315 ;
        RECT 139.090 167.085 139.550 167.315 ;
        RECT 139.880 167.085 140.340 167.315 ;
        RECT 140.670 167.085 141.130 167.315 ;
        RECT 142.920 167.085 143.380 167.315 ;
        RECT 143.710 167.085 144.170 167.315 ;
        RECT 144.500 167.085 144.960 167.315 ;
        RECT 145.290 167.085 145.750 167.315 ;
        RECT 147.540 167.085 148.000 167.315 ;
        RECT 148.330 167.085 148.790 167.315 ;
        RECT 149.120 167.085 149.580 167.315 ;
        RECT 149.910 167.085 150.370 167.315 ;
        RECT 151.150 166.625 152.755 176.325 ;
        RECT 110.685 166.035 152.755 166.625 ;
        RECT 107.745 163.060 108.705 163.290 ;
        RECT 109.035 163.060 109.995 163.290 ;
        RECT 107.745 162.990 108.445 163.060 ;
        RECT 109.295 162.990 109.995 163.060 ;
        RECT 110.685 162.685 114.420 166.035 ;
        RECT 134.745 165.030 135.445 165.080 ;
        RECT 146.905 165.030 147.605 165.080 ;
        RECT 134.745 164.430 147.605 165.030 ;
        RECT 134.745 164.380 135.445 164.430 ;
        RECT 146.905 164.380 147.605 164.430 ;
        RECT 133.735 163.740 134.435 163.790 ;
        RECT 143.985 163.740 144.685 163.790 ;
        RECT 133.735 163.140 144.685 163.740 ;
        RECT 133.735 163.090 134.435 163.140 ;
        RECT 143.985 163.090 144.685 163.140 ;
        RECT 101.935 162.285 114.420 162.685 ;
        RECT 101.935 158.755 103.025 162.285 ;
        RECT 103.435 160.445 103.665 161.520 ;
        RECT 103.400 159.745 103.700 160.445 ;
        RECT 103.435 159.520 103.665 159.745 ;
        RECT 104.725 159.520 104.955 162.285 ;
        RECT 106.015 160.445 106.245 161.520 ;
        RECT 105.980 159.745 106.280 160.445 ;
        RECT 106.015 159.520 106.245 159.745 ;
        RECT 103.715 159.130 104.675 159.360 ;
        RECT 105.005 159.130 105.965 159.360 ;
        RECT 103.845 159.060 104.545 159.130 ;
        RECT 105.135 159.060 105.835 159.130 ;
        RECT 106.655 158.755 107.055 162.285 ;
        RECT 107.465 160.445 107.695 161.520 ;
        RECT 107.430 159.745 107.730 160.445 ;
        RECT 107.465 159.520 107.695 159.745 ;
        RECT 108.755 159.520 108.985 162.285 ;
        RECT 110.045 160.445 110.275 161.520 ;
        RECT 110.010 159.745 110.310 160.445 ;
        RECT 110.045 159.520 110.275 159.745 ;
        RECT 107.745 159.130 108.705 159.360 ;
        RECT 109.035 159.130 109.995 159.360 ;
        RECT 107.875 159.060 108.575 159.130 ;
        RECT 109.165 159.060 109.865 159.130 ;
        RECT 110.685 158.755 114.420 162.285 ;
        RECT 136.825 162.330 137.525 162.400 ;
        RECT 143.985 162.330 144.685 162.400 ;
        RECT 136.825 161.730 144.685 162.330 ;
        RECT 136.825 161.700 137.525 161.730 ;
        RECT 143.985 161.700 144.685 161.730 ;
        RECT 134.745 160.160 135.445 160.210 ;
        RECT 145.575 160.160 146.275 160.210 ;
        RECT 134.745 159.560 146.275 160.160 ;
        RECT 134.745 159.510 135.445 159.560 ;
        RECT 145.575 159.510 146.275 159.560 ;
        RECT 101.935 157.850 114.420 158.755 ;
        RECT 141.665 159.150 142.365 159.200 ;
        RECT 148.605 159.150 149.305 159.200 ;
        RECT 141.665 158.550 149.305 159.150 ;
        RECT 141.665 158.500 142.365 158.550 ;
        RECT 148.605 158.500 149.305 158.550 ;
        RECT 153.960 158.060 155.900 180.110 ;
        RECT 165.150 179.490 239.210 179.970 ;
        RECT 170.755 179.290 171.045 179.335 ;
        RECT 171.200 179.290 171.520 179.350 ;
        RECT 170.755 179.150 171.520 179.290 ;
        RECT 170.755 179.105 171.045 179.150 ;
        RECT 171.200 179.090 171.520 179.150 ;
        RECT 175.340 179.090 175.660 179.350 ;
        RECT 176.260 179.290 176.580 179.350 ;
        RECT 176.735 179.290 177.025 179.335 ;
        RECT 176.260 179.150 177.025 179.290 ;
        RECT 176.260 179.090 176.580 179.150 ;
        RECT 176.735 179.105 177.025 179.150 ;
        RECT 178.560 179.290 178.880 179.350 ;
        RECT 182.715 179.290 183.005 179.335 ;
        RECT 178.560 179.150 183.005 179.290 ;
        RECT 178.560 179.090 178.880 179.150 ;
        RECT 182.715 179.105 183.005 179.150 ;
        RECT 190.060 179.290 190.380 179.350 ;
        RECT 192.835 179.290 193.125 179.335 ;
        RECT 190.060 179.150 193.125 179.290 ;
        RECT 190.060 179.090 190.380 179.150 ;
        RECT 192.835 179.105 193.125 179.150 ;
        RECT 194.200 179.290 194.520 179.350 ;
        RECT 194.200 179.150 195.810 179.290 ;
        RECT 194.200 179.090 194.520 179.150 ;
        RECT 166.600 178.950 166.920 179.010 ;
        RECT 177.640 178.950 177.960 179.010 ;
        RECT 166.600 178.810 177.960 178.950 ;
        RECT 166.600 178.750 166.920 178.810 ;
        RECT 177.640 178.750 177.960 178.810 ;
        RECT 180.875 178.950 181.165 178.995 ;
        RECT 190.535 178.950 190.825 178.995 ;
        RECT 194.660 178.950 194.980 179.010 ;
        RECT 180.875 178.810 190.295 178.950 ;
        RECT 180.875 178.765 181.165 178.810 ;
        RECT 180.400 178.610 180.720 178.670 ;
        RECT 167.150 178.470 180.720 178.610 ;
        RECT 167.150 178.315 167.290 178.470 ;
        RECT 180.400 178.410 180.720 178.470 ;
        RECT 183.710 178.470 187.990 178.610 ;
        RECT 167.075 178.085 167.365 178.315 ;
        RECT 168.440 178.070 168.760 178.330 ;
        RECT 170.740 178.315 171.060 178.330 ;
        RECT 169.835 178.085 170.125 178.315 ;
        RECT 170.605 178.270 171.060 178.315 ;
        RECT 172.120 178.270 172.440 178.330 ;
        RECT 170.605 178.130 172.440 178.270 ;
        RECT 170.605 178.085 171.060 178.130 ;
        RECT 169.910 177.930 170.050 178.085 ;
        RECT 170.740 178.070 171.060 178.085 ;
        RECT 172.120 178.070 172.440 178.130 ;
        RECT 172.580 178.270 172.900 178.330 ;
        RECT 173.055 178.270 173.345 178.315 ;
        RECT 172.580 178.130 173.345 178.270 ;
        RECT 172.580 178.070 172.900 178.130 ;
        RECT 173.055 178.085 173.345 178.130 ;
        RECT 174.420 178.070 174.740 178.330 ;
        RECT 175.815 178.085 176.105 178.315 ;
        RECT 176.280 178.085 176.570 178.315 ;
        RECT 178.575 178.085 178.865 178.315 ;
        RECT 175.890 177.930 176.030 178.085 ;
        RECT 168.070 177.790 170.050 177.930 ;
        RECT 171.810 177.790 176.030 177.930 ;
        RECT 168.070 177.635 168.210 177.790 ;
        RECT 167.995 177.405 168.285 177.635 ;
        RECT 169.375 177.590 169.665 177.635 ;
        RECT 171.810 177.590 171.950 177.790 ;
        RECT 169.375 177.450 171.950 177.590 ;
        RECT 172.120 177.590 172.440 177.650 ;
        RECT 176.350 177.590 176.490 178.085 ;
        RECT 178.650 177.930 178.790 178.085 ;
        RECT 179.940 178.070 180.260 178.330 ;
        RECT 181.320 178.070 181.640 178.330 ;
        RECT 183.710 178.315 183.850 178.470 ;
        RECT 183.635 178.085 183.925 178.315 ;
        RECT 184.095 178.270 184.385 178.315 ;
        RECT 186.380 178.270 186.700 178.330 ;
        RECT 184.095 178.130 186.700 178.270 ;
        RECT 184.095 178.085 184.385 178.130 ;
        RECT 186.380 178.070 186.700 178.130 ;
        RECT 187.300 178.070 187.620 178.330 ;
        RECT 187.850 178.270 187.990 178.470 ;
        RECT 188.220 178.410 188.540 178.670 ;
        RECT 190.155 178.610 190.295 178.810 ;
        RECT 190.535 178.810 194.980 178.950 ;
        RECT 190.535 178.765 190.825 178.810 ;
        RECT 194.660 178.750 194.980 178.810 ;
        RECT 195.670 178.655 195.810 179.150 ;
        RECT 197.880 179.090 198.200 179.350 ;
        RECT 198.355 179.290 198.645 179.335 ;
        RECT 199.260 179.290 199.580 179.350 ;
        RECT 198.355 179.150 199.580 179.290 ;
        RECT 198.355 179.105 198.645 179.150 ;
        RECT 199.260 179.090 199.580 179.150 ;
        RECT 203.400 179.090 203.720 179.350 ;
        RECT 206.620 179.290 206.940 179.350 ;
        RECT 207.095 179.290 207.385 179.335 ;
        RECT 206.620 179.150 207.385 179.290 ;
        RECT 206.620 179.090 206.940 179.150 ;
        RECT 207.095 179.105 207.385 179.150 ;
        RECT 209.380 179.290 209.700 179.350 ;
        RECT 213.520 179.290 213.840 179.350 ;
        RECT 209.380 179.150 213.840 179.290 ;
        RECT 209.380 179.090 209.700 179.150 ;
        RECT 213.150 178.995 213.290 179.150 ;
        RECT 213.520 179.090 213.840 179.150 ;
        RECT 214.900 179.290 215.220 179.350 ;
        RECT 228.240 179.290 228.560 179.350 ;
        RECT 229.175 179.290 229.465 179.335 ;
        RECT 214.900 179.150 228.010 179.290 ;
        RECT 214.900 179.090 215.220 179.150 ;
        RECT 208.885 178.950 209.175 178.995 ;
        RECT 212.115 178.950 212.405 178.995 ;
        RECT 208.885 178.810 212.405 178.950 ;
        RECT 208.885 178.765 209.175 178.810 ;
        RECT 212.115 178.765 212.405 178.810 ;
        RECT 213.075 178.765 213.365 178.995 ;
        RECT 215.820 178.750 216.140 179.010 ;
        RECT 219.515 178.950 219.805 178.995 ;
        RECT 224.155 178.950 224.445 178.995 ;
        RECT 227.385 178.950 227.675 178.995 ;
        RECT 219.515 178.810 221.110 178.950 ;
        RECT 219.515 178.765 219.805 178.810 ;
        RECT 190.155 178.470 195.350 178.610 ;
        RECT 189.615 178.270 189.905 178.315 ;
        RECT 190.980 178.270 191.300 178.330 ;
        RECT 187.850 178.130 189.370 178.270 ;
        RECT 182.700 177.930 183.020 177.990 ;
        RECT 187.775 177.930 188.065 177.975 ;
        RECT 178.650 177.790 183.020 177.930 ;
        RECT 182.700 177.730 183.020 177.790 ;
        RECT 185.090 177.790 188.065 177.930 ;
        RECT 189.230 177.930 189.370 178.130 ;
        RECT 189.615 178.130 191.300 178.270 ;
        RECT 189.615 178.085 189.905 178.130 ;
        RECT 190.980 178.070 191.300 178.130 ;
        RECT 191.455 178.270 191.745 178.315 ;
        RECT 191.900 178.270 192.220 178.330 ;
        RECT 191.455 178.130 192.220 178.270 ;
        RECT 191.455 178.085 191.745 178.130 ;
        RECT 191.900 178.070 192.220 178.130 ;
        RECT 192.820 178.270 193.140 178.330 ;
        RECT 194.675 178.270 194.965 178.315 ;
        RECT 192.820 178.130 194.965 178.270 ;
        RECT 195.210 178.270 195.350 178.470 ;
        RECT 195.595 178.425 195.885 178.655 ;
        RECT 201.100 178.610 201.420 178.670 ;
        RECT 202.020 178.610 202.340 178.670 ;
        RECT 201.100 178.470 202.340 178.610 ;
        RECT 201.100 178.410 201.420 178.470 ;
        RECT 202.020 178.410 202.340 178.470 ;
        RECT 207.540 178.610 207.860 178.670 ;
        RECT 210.300 178.610 210.620 178.670 ;
        RECT 207.540 178.470 210.620 178.610 ;
        RECT 207.540 178.410 207.860 178.470 ;
        RECT 210.300 178.410 210.620 178.470 ;
        RECT 211.110 178.610 211.400 178.655 ;
        RECT 211.110 178.470 214.670 178.610 ;
        RECT 211.110 178.425 211.400 178.470 ;
        RECT 195.210 178.130 195.810 178.270 ;
        RECT 192.820 178.070 193.140 178.130 ;
        RECT 194.675 178.085 194.965 178.130 ;
        RECT 190.060 177.930 190.380 177.990 ;
        RECT 195.135 177.930 195.425 177.975 ;
        RECT 189.230 177.790 190.380 177.930 ;
        RECT 172.120 177.450 176.490 177.590 ;
        RECT 179.495 177.590 179.785 177.635 ;
        RECT 180.860 177.590 181.180 177.650 ;
        RECT 179.495 177.450 181.180 177.590 ;
        RECT 169.375 177.405 169.665 177.450 ;
        RECT 172.120 177.390 172.440 177.450 ;
        RECT 179.495 177.405 179.785 177.450 ;
        RECT 180.860 177.390 181.180 177.450 ;
        RECT 181.780 177.590 182.100 177.650 ;
        RECT 185.090 177.635 185.230 177.790 ;
        RECT 187.775 177.745 188.065 177.790 ;
        RECT 190.060 177.730 190.380 177.790 ;
        RECT 193.370 177.790 195.425 177.930 ;
        RECT 182.255 177.590 182.545 177.635 ;
        RECT 181.780 177.450 182.545 177.590 ;
        RECT 181.780 177.390 182.100 177.450 ;
        RECT 182.255 177.405 182.545 177.450 ;
        RECT 185.015 177.405 185.305 177.635 ;
        RECT 185.475 177.590 185.765 177.635 ;
        RECT 187.300 177.590 187.620 177.650 ;
        RECT 185.475 177.450 187.620 177.590 ;
        RECT 185.475 177.405 185.765 177.450 ;
        RECT 187.300 177.390 187.620 177.450 ;
        RECT 192.375 177.590 192.665 177.635 ;
        RECT 193.370 177.590 193.510 177.790 ;
        RECT 195.135 177.745 195.425 177.790 ;
        RECT 192.375 177.450 193.510 177.590 ;
        RECT 195.670 177.590 195.810 178.130 ;
        RECT 196.975 178.085 197.265 178.315 ;
        RECT 200.655 178.270 200.945 178.315 ;
        RECT 201.560 178.270 201.880 178.330 ;
        RECT 200.655 178.130 201.880 178.270 ;
        RECT 200.655 178.085 200.945 178.130 ;
        RECT 197.050 177.930 197.190 178.085 ;
        RECT 201.560 178.070 201.880 178.130 ;
        RECT 202.495 178.270 202.785 178.315 ;
        RECT 203.400 178.270 203.720 178.330 ;
        RECT 202.495 178.130 203.720 178.270 ;
        RECT 202.495 178.085 202.785 178.130 ;
        RECT 203.400 178.070 203.720 178.130 ;
        RECT 204.320 178.270 204.640 178.330 ;
        RECT 204.795 178.270 205.085 178.315 ;
        RECT 204.320 178.130 205.085 178.270 ;
        RECT 204.320 178.070 204.640 178.130 ;
        RECT 204.795 178.085 205.085 178.130 ;
        RECT 207.965 178.270 208.255 178.315 ;
        RECT 209.805 178.270 210.095 178.315 ;
        RECT 207.965 178.130 210.095 178.270 ;
        RECT 207.965 178.085 208.255 178.130 ;
        RECT 209.805 178.085 210.095 178.130 ;
        RECT 211.680 178.070 212.000 178.330 ;
        RECT 212.150 178.270 212.440 178.315 ;
        RECT 213.990 178.270 214.280 178.315 ;
        RECT 212.150 178.130 214.280 178.270 ;
        RECT 214.530 178.270 214.670 178.470 ;
        RECT 214.900 178.410 215.220 178.670 ;
        RECT 215.910 178.610 216.050 178.750 ;
        RECT 220.970 178.655 221.110 178.810 ;
        RECT 224.155 178.810 227.675 178.950 ;
        RECT 227.870 178.950 228.010 179.150 ;
        RECT 228.240 179.150 229.465 179.290 ;
        RECT 228.240 179.090 228.560 179.150 ;
        RECT 229.175 179.105 229.465 179.150 ;
        RECT 230.095 179.290 230.385 179.335 ;
        RECT 230.540 179.290 230.860 179.350 ;
        RECT 230.095 179.150 230.860 179.290 ;
        RECT 230.095 179.105 230.385 179.150 ;
        RECT 230.540 179.090 230.860 179.150 ;
        RECT 231.460 179.090 231.780 179.350 ;
        RECT 232.380 179.290 232.700 179.350 ;
        RECT 234.235 179.290 234.525 179.335 ;
        RECT 232.380 179.150 234.525 179.290 ;
        RECT 232.380 179.090 232.700 179.150 ;
        RECT 234.235 179.105 234.525 179.150 ;
        RECT 234.680 179.290 235.000 179.350 ;
        RECT 235.615 179.290 235.905 179.335 ;
        RECT 234.680 179.150 235.905 179.290 ;
        RECT 234.680 179.090 235.000 179.150 ;
        RECT 235.615 179.105 235.905 179.150 ;
        RECT 232.855 178.950 233.145 178.995 ;
        RECT 227.870 178.810 233.145 178.950 ;
        RECT 224.155 178.765 224.445 178.810 ;
        RECT 227.385 178.765 227.675 178.810 ;
        RECT 232.855 178.765 233.145 178.810 ;
        RECT 216.295 178.610 216.585 178.655 ;
        RECT 215.910 178.470 216.585 178.610 ;
        RECT 216.295 178.425 216.585 178.470 ;
        RECT 220.895 178.425 221.185 178.655 ;
        RECT 221.340 178.610 221.660 178.670 ;
        RECT 223.195 178.610 223.485 178.655 ;
        RECT 221.340 178.470 223.485 178.610 ;
        RECT 221.340 178.410 221.660 178.470 ;
        RECT 223.195 178.425 223.485 178.470 ;
        RECT 225.265 178.610 225.555 178.655 ;
        RECT 230.080 178.610 230.400 178.670 ;
        RECT 225.265 178.470 230.400 178.610 ;
        RECT 225.265 178.425 225.555 178.470 ;
        RECT 230.080 178.410 230.400 178.470 ;
        RECT 214.990 178.270 215.130 178.410 ;
        RECT 214.530 178.130 215.130 178.270 ;
        RECT 212.150 178.085 212.440 178.130 ;
        RECT 213.990 178.085 214.280 178.130 ;
        RECT 215.375 178.085 215.665 178.315 ;
        RECT 215.820 178.270 216.140 178.330 ;
        RECT 217.215 178.270 217.505 178.315 ;
        RECT 215.820 178.130 217.505 178.270 ;
        RECT 208.470 177.930 208.760 177.975 ;
        RECT 209.390 177.930 209.680 177.975 ;
        RECT 214.910 177.930 215.200 177.975 ;
        RECT 197.050 177.790 201.790 177.930 ;
        RECT 201.650 177.650 201.790 177.790 ;
        RECT 208.470 177.790 215.200 177.930 ;
        RECT 208.470 177.745 208.760 177.790 ;
        RECT 209.390 177.745 209.680 177.790 ;
        RECT 214.910 177.745 215.200 177.790 ;
        RECT 200.195 177.590 200.485 177.635 ;
        RECT 195.670 177.450 200.485 177.590 ;
        RECT 192.375 177.405 192.665 177.450 ;
        RECT 200.195 177.405 200.485 177.450 ;
        RECT 201.560 177.390 201.880 177.650 ;
        RECT 205.715 177.590 206.005 177.635 ;
        RECT 215.450 177.590 215.590 178.085 ;
        RECT 215.820 178.070 216.140 178.130 ;
        RECT 217.215 178.085 217.505 178.130 ;
        RECT 217.660 178.270 217.980 178.330 ;
        RECT 218.595 178.270 218.885 178.315 ;
        RECT 217.660 178.130 218.885 178.270 ;
        RECT 217.660 178.070 217.980 178.130 ;
        RECT 218.595 178.085 218.885 178.130 ;
        RECT 219.500 178.270 219.820 178.330 ;
        RECT 219.975 178.270 220.265 178.315 ;
        RECT 219.500 178.130 220.265 178.270 ;
        RECT 219.500 178.070 219.820 178.130 ;
        RECT 219.975 178.085 220.265 178.130 ;
        RECT 222.280 178.270 222.570 178.315 ;
        RECT 224.120 178.270 224.410 178.315 ;
        RECT 222.280 178.130 224.410 178.270 ;
        RECT 222.280 178.085 222.570 178.130 ;
        RECT 224.120 178.085 224.410 178.130 ;
        RECT 224.560 178.070 224.880 178.330 ;
        RECT 225.940 178.070 226.260 178.330 ;
        RECT 226.465 178.270 226.755 178.315 ;
        RECT 228.305 178.270 228.595 178.315 ;
        RECT 226.465 178.130 228.595 178.270 ;
        RECT 226.465 178.085 226.755 178.130 ;
        RECT 228.305 178.085 228.595 178.130 ;
        RECT 229.620 178.270 229.940 178.330 ;
        RECT 231.015 178.270 231.305 178.315 ;
        RECT 229.620 178.130 231.305 178.270 ;
        RECT 229.620 178.070 229.940 178.130 ;
        RECT 231.015 178.085 231.305 178.130 ;
        RECT 232.380 178.070 232.700 178.330 ;
        RECT 233.760 178.070 234.080 178.330 ;
        RECT 235.155 178.085 235.445 178.315 ;
        RECT 221.360 177.930 221.650 177.975 ;
        RECT 226.880 177.930 227.170 177.975 ;
        RECT 227.800 177.930 228.090 177.975 ;
        RECT 235.230 177.930 235.370 178.085 ;
        RECT 236.520 178.070 236.840 178.330 ;
        RECT 221.360 177.790 228.090 177.930 ;
        RECT 221.360 177.745 221.650 177.790 ;
        RECT 226.880 177.745 227.170 177.790 ;
        RECT 227.800 177.745 228.090 177.790 ;
        RECT 229.710 177.790 235.370 177.930 ;
        RECT 205.715 177.450 215.590 177.590 ;
        RECT 218.135 177.590 218.425 177.635 ;
        RECT 220.420 177.590 220.740 177.650 ;
        RECT 218.135 177.450 220.740 177.590 ;
        RECT 205.715 177.405 206.005 177.450 ;
        RECT 218.135 177.405 218.425 177.450 ;
        RECT 220.420 177.390 220.740 177.450 ;
        RECT 220.880 177.590 221.200 177.650 ;
        RECT 229.710 177.590 229.850 177.790 ;
        RECT 220.880 177.450 229.850 177.590 ;
        RECT 220.880 177.390 221.200 177.450 ;
        RECT 165.150 176.770 239.210 177.250 ;
        RECT 185.460 176.370 185.780 176.630 ;
        RECT 191.900 176.570 192.220 176.630 ;
        RECT 198.340 176.570 198.660 176.630 ;
        RECT 191.900 176.430 198.660 176.570 ;
        RECT 191.900 176.370 192.220 176.430 ;
        RECT 198.340 176.370 198.660 176.430 ;
        RECT 207.540 176.570 207.860 176.630 ;
        RECT 215.820 176.570 216.140 176.630 ;
        RECT 207.540 176.430 216.140 176.570 ;
        RECT 207.540 176.370 207.860 176.430 ;
        RECT 215.820 176.370 216.140 176.430 ;
        RECT 225.940 176.570 226.260 176.630 ;
        RECT 235.140 176.570 235.460 176.630 ;
        RECT 225.940 176.430 235.460 176.570 ;
        RECT 225.940 176.370 226.260 176.430 ;
        RECT 235.140 176.370 235.460 176.430 ;
        RECT 177.180 176.230 177.500 176.290 ;
        RECT 185.550 176.230 185.690 176.370 ;
        RECT 187.300 176.230 187.620 176.290 ;
        RECT 177.180 176.090 185.690 176.230 ;
        RECT 186.010 176.090 187.620 176.230 ;
        RECT 177.180 176.030 177.500 176.090 ;
        RECT 178.100 175.890 178.420 175.950 ;
        RECT 186.010 175.890 186.150 176.090 ;
        RECT 187.300 176.030 187.620 176.090 ;
        RECT 208.460 176.230 208.780 176.290 ;
        RECT 217.660 176.230 217.980 176.290 ;
        RECT 221.340 176.230 221.660 176.290 ;
        RECT 208.460 176.090 217.980 176.230 ;
        RECT 208.460 176.030 208.780 176.090 ;
        RECT 217.660 176.030 217.980 176.090 ;
        RECT 219.130 176.090 221.660 176.230 ;
        RECT 178.100 175.750 186.150 175.890 ;
        RECT 186.380 175.890 186.700 175.950 ;
        RECT 195.580 175.890 195.900 175.950 ;
        RECT 186.380 175.750 195.900 175.890 ;
        RECT 178.100 175.690 178.420 175.750 ;
        RECT 186.380 175.690 186.700 175.750 ;
        RECT 195.580 175.690 195.900 175.750 ;
        RECT 202.020 175.890 202.340 175.950 ;
        RECT 219.130 175.890 219.270 176.090 ;
        RECT 221.340 176.030 221.660 176.090 ;
        RECT 222.260 176.230 222.580 176.290 ;
        RECT 236.520 176.230 236.840 176.290 ;
        RECT 222.260 176.090 236.840 176.230 ;
        RECT 222.260 176.030 222.580 176.090 ;
        RECT 236.520 176.030 236.840 176.090 ;
        RECT 202.020 175.750 219.270 175.890 ;
        RECT 219.500 175.890 219.820 175.950 ;
        RECT 233.760 175.890 234.080 175.950 ;
        RECT 219.500 175.750 234.080 175.890 ;
        RECT 202.020 175.690 202.340 175.750 ;
        RECT 219.500 175.690 219.820 175.750 ;
        RECT 233.760 175.690 234.080 175.750 ;
        RECT 179.940 175.550 180.260 175.610 ;
        RECT 192.820 175.550 193.140 175.610 ;
        RECT 179.940 175.410 193.140 175.550 ;
        RECT 179.940 175.350 180.260 175.410 ;
        RECT 192.820 175.350 193.140 175.410 ;
        RECT 218.580 175.550 218.900 175.610 ;
        RECT 232.380 175.550 232.700 175.610 ;
        RECT 218.580 175.410 232.700 175.550 ;
        RECT 218.580 175.350 218.900 175.410 ;
        RECT 232.380 175.350 232.700 175.410 ;
        RECT 181.780 175.210 182.100 175.270 ;
        RECT 196.500 175.210 196.820 175.270 ;
        RECT 181.780 175.070 196.820 175.210 ;
        RECT 181.780 175.010 182.100 175.070 ;
        RECT 196.500 175.010 196.820 175.070 ;
        RECT 216.740 175.210 217.060 175.270 ;
        RECT 229.620 175.210 229.940 175.270 ;
        RECT 216.740 175.070 229.940 175.210 ;
        RECT 216.740 175.010 217.060 175.070 ;
        RECT 229.620 175.010 229.940 175.070 ;
        RECT 180.860 174.870 181.180 174.930 ;
        RECT 193.740 174.870 194.060 174.930 ;
        RECT 180.860 174.730 194.060 174.870 ;
        RECT 180.860 174.670 181.180 174.730 ;
        RECT 193.740 174.670 194.060 174.730 ;
        RECT 190.060 174.530 190.380 174.590 ;
        RECT 194.660 174.530 194.980 174.590 ;
        RECT 190.060 174.390 194.980 174.530 ;
        RECT 190.060 174.330 190.380 174.390 ;
        RECT 194.660 174.330 194.980 174.390 ;
        RECT 115.985 156.185 155.900 158.060 ;
        RECT 115.985 156.060 116.575 156.185 ;
        RECT 102.625 155.660 116.575 156.060 ;
        RECT 102.625 152.040 103.025 155.660 ;
        RECT 103.715 155.055 104.675 155.385 ;
        RECT 105.005 155.055 105.965 155.385 ;
        RECT 103.435 153.515 103.665 154.850 ;
        RECT 103.400 152.815 103.700 153.515 ;
        RECT 104.725 152.040 104.955 154.850 ;
        RECT 106.015 154.585 106.245 154.850 ;
        RECT 105.980 153.885 106.280 154.585 ;
        RECT 106.015 152.850 106.245 153.885 ;
        RECT 106.655 152.040 107.055 155.660 ;
        RECT 107.745 155.055 108.705 155.385 ;
        RECT 109.035 155.055 109.995 155.385 ;
        RECT 107.465 153.515 107.695 154.850 ;
        RECT 107.430 152.815 107.730 153.515 ;
        RECT 108.755 152.040 108.985 154.850 ;
        RECT 110.045 154.585 110.275 154.850 ;
        RECT 110.010 153.885 110.310 154.585 ;
        RECT 110.045 152.850 110.275 153.885 ;
        RECT 110.685 152.040 116.575 155.660 ;
        RECT 102.625 151.550 116.575 152.040 ;
        RECT 102.625 142.020 103.025 151.550 ;
        RECT 103.715 151.035 104.675 151.365 ;
        RECT 105.005 151.035 105.965 151.365 ;
        RECT 103.435 145.785 103.665 150.830 ;
        RECT 104.725 149.485 104.955 150.830 ;
        RECT 104.690 147.185 104.990 149.485 ;
        RECT 103.400 143.485 103.700 145.785 ;
        RECT 103.435 142.830 103.665 143.485 ;
        RECT 104.725 142.830 104.955 147.185 ;
        RECT 106.015 145.785 106.245 150.830 ;
        RECT 105.980 143.485 106.280 145.785 ;
        RECT 106.015 142.830 106.245 143.485 ;
        RECT 103.715 142.395 104.675 142.625 ;
        RECT 105.005 142.395 105.965 142.625 ;
        RECT 106.655 142.020 107.055 151.550 ;
        RECT 107.745 151.035 108.705 151.365 ;
        RECT 109.035 151.035 109.995 151.365 ;
        RECT 107.465 145.785 107.695 150.830 ;
        RECT 108.755 149.485 108.985 150.830 ;
        RECT 108.720 147.185 109.020 149.485 ;
        RECT 107.430 143.485 107.730 145.785 ;
        RECT 107.465 142.830 107.695 143.485 ;
        RECT 108.755 142.830 108.985 147.185 ;
        RECT 110.045 145.785 110.275 150.830 ;
        RECT 110.010 143.485 110.310 145.785 ;
        RECT 110.045 142.830 110.275 143.485 ;
        RECT 107.745 142.395 108.705 142.625 ;
        RECT 109.035 142.395 109.995 142.625 ;
        RECT 110.685 142.020 116.575 151.550 ;
        RECT 117.160 142.145 119.265 155.605 ;
        RECT 122.405 146.245 124.510 155.605 ;
        RECT 125.090 146.825 127.195 155.605 ;
        RECT 130.335 146.825 132.440 155.605 ;
        RECT 133.020 154.960 135.125 155.660 ;
        RECT 133.020 152.675 135.125 154.435 ;
        RECT 138.265 153.845 140.370 155.605 ;
        RECT 133.020 151.450 135.125 152.150 ;
        RECT 138.265 151.505 140.370 153.265 ;
        RECT 140.950 152.675 143.055 156.185 ;
        RECT 146.195 152.675 148.300 156.185 ;
        RECT 140.950 151.460 143.055 152.160 ;
        RECT 133.020 150.280 135.125 150.980 ;
        RECT 133.020 149.110 135.125 149.810 ;
        RECT 138.265 149.165 140.370 150.925 ;
        RECT 140.950 149.165 143.055 150.925 ;
        RECT 146.195 150.335 148.300 152.095 ;
        RECT 133.020 146.825 135.125 148.585 ;
        RECT 138.265 146.825 140.370 148.585 ;
        RECT 140.950 146.825 143.055 148.585 ;
        RECT 146.195 147.995 148.300 149.755 ;
        RECT 122.405 142.145 127.195 146.245 ;
        RECT 130.335 142.145 132.440 146.245 ;
        RECT 133.020 142.145 135.125 146.245 ;
        RECT 138.265 142.145 140.370 146.245 ;
        RECT 140.950 144.485 143.055 146.245 ;
        RECT 146.195 145.655 148.300 147.415 ;
        RECT 140.950 143.290 143.055 143.990 ;
        RECT 146.195 143.315 148.300 145.075 ;
        RECT 140.950 142.040 143.055 142.740 ;
        RECT 146.195 142.080 148.300 142.780 ;
        RECT 102.625 141.620 116.575 142.020 ;
        RECT 62.865 130.990 100.480 139.455 ;
        RECT 111.085 141.565 116.575 141.620 ;
        RECT 148.885 141.565 155.900 156.185 ;
        RECT 111.085 137.690 155.900 141.565 ;
        RECT 111.085 130.990 135.120 137.690 ;
        RECT 62.865 127.485 135.120 130.990 ;
        RECT 138.080 134.100 145.960 137.690 ;
        RECT 138.080 130.310 138.670 134.100 ;
        RECT 139.615 133.640 140.315 133.760 ;
        RECT 140.905 133.640 141.605 133.760 ;
        RECT 139.485 133.410 140.445 133.640 ;
        RECT 140.775 133.410 141.735 133.640 ;
        RECT 139.205 132.990 139.435 133.205 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 139.205 131.205 139.435 131.390 ;
        RECT 140.495 130.310 140.725 133.205 ;
        RECT 141.785 132.990 142.015 133.205 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 143.315 132.640 143.545 133.205 ;
        RECT 143.280 131.940 143.580 132.640 ;
        RECT 141.785 131.205 142.015 131.390 ;
        RECT 143.315 131.205 143.545 131.940 ;
        RECT 144.605 131.205 144.835 134.100 ;
        RECT 143.595 130.770 144.555 131.000 ;
        RECT 143.725 130.700 144.425 130.770 ;
        RECT 145.370 130.310 145.960 134.100 ;
        RECT 138.080 129.720 145.960 130.310 ;
        RECT 4.100 124.285 135.120 127.485 ;
        RECT 4.100 44.835 4.900 124.285 ;
        RECT 8.665 123.695 70.175 124.285 ;
        RECT 8.665 122.800 10.615 123.695 ;
        RECT 11.335 123.005 13.295 123.235 ;
        RECT 13.625 123.005 15.585 123.235 ;
        RECT 17.255 123.005 19.215 123.305 ;
        RECT 19.545 123.005 21.505 123.305 ;
        RECT 23.175 123.005 25.135 123.305 ;
        RECT 25.465 123.005 27.425 123.305 ;
        RECT 29.095 123.005 31.055 123.305 ;
        RECT 31.385 123.005 33.345 123.305 ;
        RECT 35.015 123.005 36.975 123.305 ;
        RECT 37.305 123.005 39.265 123.305 ;
        RECT 40.935 123.005 42.895 123.305 ;
        RECT 43.225 123.005 45.185 123.305 ;
        RECT 46.855 123.005 48.815 123.305 ;
        RECT 49.145 123.005 51.105 123.305 ;
        RECT 52.775 123.005 54.735 123.305 ;
        RECT 55.065 123.005 57.025 123.305 ;
        RECT 58.695 123.005 60.655 123.305 ;
        RECT 60.985 123.005 62.945 123.305 ;
        RECT 64.615 123.005 66.575 123.235 ;
        RECT 66.905 123.005 68.865 123.235 ;
        RECT 69.585 122.800 70.175 123.695 ;
        RECT 8.665 117.050 11.285 122.800 ;
        RECT 13.345 117.050 13.575 122.800 ;
        RECT 15.635 117.050 15.865 122.800 ;
        RECT 16.975 117.050 17.205 122.800 ;
        RECT 19.265 122.050 19.495 122.800 ;
        RECT 19.030 120.550 19.730 122.050 ;
        RECT 8.665 115.550 11.520 117.050 ;
        RECT 13.110 115.550 13.810 117.050 ;
        RECT 15.400 115.550 16.100 117.050 ;
        RECT 16.740 115.550 17.440 117.050 ;
        RECT 8.665 114.595 11.285 115.550 ;
        RECT 13.345 114.595 13.575 115.550 ;
        RECT 15.635 114.595 15.865 115.550 ;
        RECT 16.975 114.800 17.205 115.550 ;
        RECT 19.265 114.800 19.495 120.550 ;
        RECT 21.555 117.050 21.785 122.800 ;
        RECT 22.895 117.050 23.125 122.800 ;
        RECT 25.185 119.550 25.415 122.800 ;
        RECT 24.950 118.050 25.650 119.550 ;
        RECT 21.320 115.550 22.020 117.050 ;
        RECT 22.660 115.550 23.360 117.050 ;
        RECT 21.555 114.800 21.785 115.550 ;
        RECT 22.895 114.800 23.125 115.550 ;
        RECT 25.185 114.800 25.415 118.050 ;
        RECT 27.475 117.050 27.705 122.800 ;
        RECT 28.815 117.050 29.045 122.800 ;
        RECT 27.240 115.550 27.940 117.050 ;
        RECT 28.580 115.550 29.280 117.050 ;
        RECT 27.475 114.800 27.705 115.550 ;
        RECT 28.815 114.800 29.045 115.550 ;
        RECT 31.105 114.595 31.335 122.800 ;
        RECT 33.395 117.050 33.625 122.800 ;
        RECT 34.735 117.050 34.965 122.800 ;
        RECT 37.025 122.050 37.255 122.800 ;
        RECT 36.790 120.550 37.490 122.050 ;
        RECT 33.160 115.550 33.860 117.050 ;
        RECT 34.500 115.550 35.200 117.050 ;
        RECT 33.395 114.800 33.625 115.550 ;
        RECT 34.735 114.800 34.965 115.550 ;
        RECT 37.025 114.800 37.255 120.550 ;
        RECT 39.315 117.050 39.545 122.800 ;
        RECT 40.655 117.050 40.885 122.800 ;
        RECT 42.945 122.050 43.175 122.800 ;
        RECT 42.710 120.550 43.410 122.050 ;
        RECT 39.080 115.550 39.780 117.050 ;
        RECT 40.420 115.550 41.120 117.050 ;
        RECT 39.315 114.800 39.545 115.550 ;
        RECT 40.655 114.800 40.885 115.550 ;
        RECT 42.945 114.800 43.175 120.550 ;
        RECT 45.235 117.050 45.465 122.800 ;
        RECT 46.575 117.050 46.805 122.800 ;
        RECT 45.000 115.550 45.700 117.050 ;
        RECT 46.340 115.550 47.040 117.050 ;
        RECT 45.235 114.800 45.465 115.550 ;
        RECT 46.575 114.800 46.805 115.550 ;
        RECT 48.865 114.595 49.095 122.800 ;
        RECT 51.155 117.050 51.385 122.800 ;
        RECT 52.495 117.050 52.725 122.800 ;
        RECT 54.785 119.550 55.015 122.800 ;
        RECT 54.550 118.050 55.250 119.550 ;
        RECT 50.920 115.550 51.620 117.050 ;
        RECT 52.260 115.550 52.960 117.050 ;
        RECT 51.155 114.800 51.385 115.550 ;
        RECT 52.495 114.800 52.725 115.550 ;
        RECT 54.785 114.800 55.015 118.050 ;
        RECT 57.075 117.050 57.305 122.800 ;
        RECT 58.415 117.050 58.645 122.800 ;
        RECT 60.705 122.050 60.935 122.800 ;
        RECT 60.470 120.550 61.170 122.050 ;
        RECT 56.840 115.550 57.540 117.050 ;
        RECT 58.180 115.550 58.880 117.050 ;
        RECT 57.075 114.800 57.305 115.550 ;
        RECT 58.415 114.800 58.645 115.550 ;
        RECT 60.705 114.800 60.935 120.550 ;
        RECT 62.995 117.050 63.225 122.800 ;
        RECT 64.335 117.050 64.565 122.800 ;
        RECT 66.625 117.050 66.855 122.800 ;
        RECT 68.915 117.050 70.175 122.800 ;
        RECT 62.760 115.550 63.460 117.050 ;
        RECT 64.100 115.550 64.800 117.050 ;
        RECT 66.390 115.550 67.090 117.050 ;
        RECT 68.680 115.550 70.175 117.050 ;
        RECT 62.995 114.800 63.225 115.550 ;
        RECT 64.335 114.595 64.565 115.550 ;
        RECT 66.625 114.595 66.855 115.550 ;
        RECT 68.915 114.595 70.175 115.550 ;
        RECT 8.665 114.365 15.865 114.595 ;
        RECT 8.665 113.215 10.615 114.365 ;
        RECT 17.255 114.295 19.215 114.595 ;
        RECT 19.545 114.295 21.505 114.595 ;
        RECT 23.175 114.295 25.135 114.595 ;
        RECT 25.465 114.295 27.425 114.595 ;
        RECT 29.095 114.365 33.345 114.595 ;
        RECT 29.095 114.295 31.055 114.365 ;
        RECT 31.385 114.295 33.345 114.365 ;
        RECT 35.015 114.295 36.975 114.595 ;
        RECT 37.305 114.295 39.265 114.595 ;
        RECT 40.935 114.295 42.895 114.595 ;
        RECT 43.225 114.295 45.185 114.595 ;
        RECT 46.855 114.365 51.105 114.595 ;
        RECT 46.855 114.295 48.815 114.365 ;
        RECT 49.145 114.295 51.105 114.365 ;
        RECT 52.775 114.295 54.735 114.595 ;
        RECT 55.065 114.295 57.025 114.595 ;
        RECT 58.695 114.295 60.655 114.595 ;
        RECT 60.985 114.295 62.945 114.595 ;
        RECT 64.335 114.365 70.175 114.595 ;
        RECT 8.665 112.985 15.865 113.215 ;
        RECT 17.255 112.985 19.215 113.285 ;
        RECT 19.545 112.985 21.505 113.285 ;
        RECT 23.175 112.985 25.135 113.285 ;
        RECT 25.465 112.985 27.425 113.285 ;
        RECT 29.095 113.215 31.055 113.285 ;
        RECT 31.385 113.215 33.345 113.285 ;
        RECT 29.095 112.985 33.345 113.215 ;
        RECT 35.015 112.985 36.975 113.285 ;
        RECT 37.305 112.985 39.265 113.285 ;
        RECT 40.935 112.985 42.895 113.285 ;
        RECT 43.225 112.985 45.185 113.285 ;
        RECT 46.855 113.215 48.815 113.285 ;
        RECT 49.145 113.215 51.105 113.285 ;
        RECT 46.855 112.985 51.105 113.215 ;
        RECT 52.775 112.985 54.735 113.285 ;
        RECT 55.065 112.985 57.025 113.285 ;
        RECT 58.695 112.985 60.655 113.285 ;
        RECT 60.985 112.985 62.945 113.285 ;
        RECT 69.585 113.215 70.175 114.365 ;
        RECT 64.335 112.985 70.175 113.215 ;
        RECT 8.665 112.030 11.285 112.985 ;
        RECT 13.345 112.030 13.575 112.985 ;
        RECT 15.635 112.030 15.865 112.985 ;
        RECT 16.975 112.030 17.205 112.780 ;
        RECT 8.665 110.530 11.520 112.030 ;
        RECT 13.110 110.530 13.810 112.030 ;
        RECT 15.400 110.530 16.100 112.030 ;
        RECT 16.740 110.530 17.440 112.030 ;
        RECT 8.665 104.780 11.285 110.530 ;
        RECT 13.345 104.780 13.575 110.530 ;
        RECT 15.635 104.780 15.865 110.530 ;
        RECT 16.975 104.780 17.205 110.530 ;
        RECT 19.265 107.030 19.495 112.780 ;
        RECT 21.555 112.030 21.785 112.780 ;
        RECT 22.895 112.030 23.125 112.780 ;
        RECT 21.320 110.530 22.020 112.030 ;
        RECT 22.660 110.530 23.360 112.030 ;
        RECT 19.030 105.530 19.730 107.030 ;
        RECT 19.265 104.780 19.495 105.530 ;
        RECT 21.555 104.780 21.785 110.530 ;
        RECT 22.895 104.780 23.125 110.530 ;
        RECT 25.185 109.530 25.415 112.780 ;
        RECT 27.475 112.030 27.705 112.780 ;
        RECT 28.815 112.030 29.045 112.780 ;
        RECT 27.240 110.530 27.940 112.030 ;
        RECT 28.580 110.530 29.280 112.030 ;
        RECT 24.950 108.030 25.650 109.530 ;
        RECT 25.185 104.780 25.415 108.030 ;
        RECT 27.475 104.780 27.705 110.530 ;
        RECT 28.815 104.780 29.045 110.530 ;
        RECT 31.105 104.780 31.335 112.985 ;
        RECT 33.395 112.030 33.625 112.780 ;
        RECT 34.735 112.030 34.965 112.780 ;
        RECT 33.160 110.530 33.860 112.030 ;
        RECT 34.500 110.530 35.200 112.030 ;
        RECT 33.395 104.780 33.625 110.530 ;
        RECT 34.735 104.780 34.965 110.530 ;
        RECT 37.025 107.030 37.255 112.780 ;
        RECT 39.315 112.030 39.545 112.780 ;
        RECT 40.655 112.030 40.885 112.780 ;
        RECT 39.080 110.530 39.780 112.030 ;
        RECT 40.420 110.530 41.120 112.030 ;
        RECT 36.790 105.530 37.490 107.030 ;
        RECT 37.025 104.780 37.255 105.530 ;
        RECT 39.315 104.780 39.545 110.530 ;
        RECT 40.655 104.780 40.885 110.530 ;
        RECT 42.945 107.030 43.175 112.780 ;
        RECT 45.235 112.030 45.465 112.780 ;
        RECT 46.575 112.030 46.805 112.780 ;
        RECT 45.000 110.530 45.700 112.030 ;
        RECT 46.340 110.530 47.040 112.030 ;
        RECT 42.710 105.530 43.410 107.030 ;
        RECT 42.945 104.780 43.175 105.530 ;
        RECT 45.235 104.780 45.465 110.530 ;
        RECT 46.575 104.780 46.805 110.530 ;
        RECT 48.865 104.780 49.095 112.985 ;
        RECT 51.155 112.030 51.385 112.780 ;
        RECT 52.495 112.030 52.725 112.780 ;
        RECT 50.920 110.530 51.620 112.030 ;
        RECT 52.260 110.530 52.960 112.030 ;
        RECT 51.155 104.780 51.385 110.530 ;
        RECT 52.495 104.780 52.725 110.530 ;
        RECT 54.785 109.530 55.015 112.780 ;
        RECT 57.075 112.030 57.305 112.780 ;
        RECT 58.415 112.030 58.645 112.780 ;
        RECT 56.840 110.530 57.540 112.030 ;
        RECT 58.180 110.530 58.880 112.030 ;
        RECT 54.550 108.030 55.250 109.530 ;
        RECT 54.785 104.780 55.015 108.030 ;
        RECT 57.075 104.780 57.305 110.530 ;
        RECT 58.415 104.780 58.645 110.530 ;
        RECT 60.705 107.030 60.935 112.780 ;
        RECT 62.995 112.030 63.225 112.780 ;
        RECT 64.335 112.030 64.565 112.985 ;
        RECT 66.625 112.030 66.855 112.985 ;
        RECT 68.915 112.030 70.175 112.985 ;
        RECT 62.760 110.530 63.460 112.030 ;
        RECT 64.100 110.530 64.800 112.030 ;
        RECT 66.390 110.530 67.090 112.030 ;
        RECT 68.680 110.530 70.175 112.030 ;
        RECT 60.470 105.530 61.170 107.030 ;
        RECT 60.705 104.780 60.935 105.530 ;
        RECT 62.995 104.780 63.225 110.530 ;
        RECT 64.335 104.780 64.565 110.530 ;
        RECT 66.625 104.780 66.855 110.530 ;
        RECT 68.915 104.780 70.175 110.530 ;
        RECT 8.665 103.885 10.615 104.780 ;
        RECT 11.335 104.345 13.295 104.575 ;
        RECT 13.625 104.345 15.585 104.575 ;
        RECT 17.255 104.275 19.215 104.575 ;
        RECT 19.545 104.275 21.505 104.575 ;
        RECT 23.175 104.275 25.135 104.575 ;
        RECT 25.465 104.275 27.425 104.575 ;
        RECT 29.095 104.275 31.055 104.575 ;
        RECT 31.385 104.275 33.345 104.575 ;
        RECT 35.015 104.275 36.975 104.575 ;
        RECT 37.305 104.275 39.265 104.575 ;
        RECT 40.935 104.275 42.895 104.575 ;
        RECT 43.225 104.275 45.185 104.575 ;
        RECT 46.855 104.275 48.815 104.575 ;
        RECT 49.145 104.275 51.105 104.575 ;
        RECT 52.775 104.275 54.735 104.575 ;
        RECT 55.065 104.275 57.025 104.575 ;
        RECT 58.695 104.275 60.655 104.575 ;
        RECT 60.985 104.275 62.945 104.575 ;
        RECT 64.615 104.345 66.575 104.575 ;
        RECT 66.905 104.345 68.865 104.575 ;
        RECT 69.585 103.885 70.175 104.780 ;
        RECT 8.665 102.705 70.175 103.885 ;
        RECT 71.775 123.695 114.165 124.285 ;
        RECT 71.775 103.885 72.365 123.695 ;
        RECT 72.805 122.800 77.615 123.695 ;
        RECT 79.005 123.005 80.965 123.305 ;
        RECT 81.295 123.005 83.255 123.305 ;
        RECT 84.925 123.005 86.885 123.305 ;
        RECT 87.215 123.005 89.175 123.305 ;
        RECT 90.845 123.005 95.095 123.305 ;
        RECT 96.765 123.005 98.725 123.305 ;
        RECT 99.055 123.005 101.015 123.305 ;
        RECT 102.685 123.005 104.645 123.305 ;
        RECT 104.975 123.005 106.935 123.305 ;
        RECT 72.805 114.800 73.035 122.800 ;
        RECT 75.095 114.800 75.325 122.800 ;
        RECT 77.385 114.800 77.615 122.800 ;
        RECT 78.725 120.650 78.955 122.800 ;
        RECT 78.490 119.950 79.190 120.650 ;
        RECT 78.725 114.800 78.955 119.950 ;
        RECT 81.015 119.150 81.245 122.800 ;
        RECT 83.305 120.650 83.535 122.800 ;
        RECT 83.070 119.950 83.770 120.650 ;
        RECT 80.780 118.450 81.480 119.150 ;
        RECT 81.015 114.800 81.245 118.450 ;
        RECT 83.305 114.800 83.535 119.950 ;
        RECT 84.645 116.150 84.875 122.800 ;
        RECT 86.935 117.650 87.165 122.800 ;
        RECT 86.700 116.950 87.400 117.650 ;
        RECT 84.410 115.450 85.110 116.150 ;
        RECT 84.645 114.800 84.875 115.450 ;
        RECT 86.935 114.800 87.165 116.950 ;
        RECT 89.225 116.150 89.455 122.800 ;
        RECT 90.565 122.150 90.795 122.800 ;
        RECT 90.330 121.450 91.030 122.150 ;
        RECT 88.990 115.450 89.690 116.150 ;
        RECT 89.225 114.800 89.455 115.450 ;
        RECT 90.565 114.800 90.795 121.450 ;
        RECT 92.855 114.800 93.085 123.005 ;
        RECT 108.325 122.800 113.135 123.695 ;
        RECT 95.145 122.150 95.375 122.800 ;
        RECT 94.910 121.450 95.610 122.150 ;
        RECT 95.145 114.800 95.375 121.450 ;
        RECT 96.485 116.150 96.715 122.800 ;
        RECT 98.775 117.650 99.005 122.800 ;
        RECT 98.540 116.950 99.240 117.650 ;
        RECT 96.250 115.450 96.950 116.150 ;
        RECT 96.485 114.800 96.715 115.450 ;
        RECT 98.775 114.800 99.005 116.950 ;
        RECT 101.065 116.150 101.295 122.800 ;
        RECT 102.405 120.650 102.635 122.800 ;
        RECT 102.170 119.950 102.870 120.650 ;
        RECT 100.830 115.450 101.530 116.150 ;
        RECT 101.065 114.800 101.295 115.450 ;
        RECT 102.405 114.800 102.635 119.950 ;
        RECT 104.695 119.150 104.925 122.800 ;
        RECT 106.985 120.650 107.215 122.800 ;
        RECT 106.750 119.950 107.450 120.650 ;
        RECT 104.460 118.450 105.160 119.150 ;
        RECT 104.695 114.800 104.925 118.450 ;
        RECT 106.985 114.800 107.215 119.950 ;
        RECT 108.325 114.800 108.555 122.800 ;
        RECT 110.615 114.800 110.845 122.800 ;
        RECT 112.905 114.800 113.135 122.800 ;
        RECT 73.085 114.365 75.045 114.595 ;
        RECT 75.375 114.365 77.335 114.595 ;
        RECT 79.005 114.295 80.965 114.595 ;
        RECT 81.295 114.295 83.255 114.595 ;
        RECT 84.925 114.295 86.885 114.595 ;
        RECT 87.215 114.295 89.175 114.595 ;
        RECT 90.845 114.295 92.805 114.595 ;
        RECT 93.135 114.295 95.095 114.595 ;
        RECT 96.765 114.295 98.725 114.595 ;
        RECT 99.055 114.295 101.015 114.595 ;
        RECT 102.685 114.295 104.645 114.595 ;
        RECT 104.975 114.295 106.935 114.595 ;
        RECT 108.605 114.365 110.565 114.595 ;
        RECT 110.895 114.365 112.855 114.595 ;
        RECT 73.085 112.985 75.045 113.215 ;
        RECT 75.375 112.985 77.335 113.215 ;
        RECT 79.005 112.985 80.965 113.285 ;
        RECT 81.295 112.985 83.255 113.285 ;
        RECT 84.925 112.985 86.885 113.285 ;
        RECT 87.215 112.985 89.175 113.285 ;
        RECT 90.845 112.985 92.805 113.285 ;
        RECT 93.135 112.985 95.095 113.285 ;
        RECT 96.765 112.985 98.725 113.285 ;
        RECT 99.055 112.985 101.015 113.285 ;
        RECT 102.685 112.985 104.645 113.285 ;
        RECT 104.975 112.985 106.935 113.285 ;
        RECT 108.605 112.985 110.565 113.215 ;
        RECT 110.895 112.985 112.855 113.215 ;
        RECT 72.805 104.780 73.035 112.780 ;
        RECT 75.095 104.780 75.325 112.780 ;
        RECT 77.385 104.780 77.615 112.780 ;
        RECT 78.725 107.630 78.955 112.780 ;
        RECT 81.015 109.130 81.245 112.780 ;
        RECT 80.780 108.430 81.480 109.130 ;
        RECT 78.490 106.930 79.190 107.630 ;
        RECT 78.725 104.780 78.955 106.930 ;
        RECT 81.015 104.780 81.245 108.430 ;
        RECT 83.305 107.630 83.535 112.780 ;
        RECT 84.645 112.130 84.875 112.780 ;
        RECT 84.410 111.430 85.110 112.130 ;
        RECT 83.070 106.930 83.770 107.630 ;
        RECT 83.305 104.780 83.535 106.930 ;
        RECT 84.645 104.780 84.875 111.430 ;
        RECT 86.935 110.630 87.165 112.780 ;
        RECT 89.225 112.130 89.455 112.780 ;
        RECT 88.990 111.430 89.690 112.130 ;
        RECT 86.700 109.930 87.400 110.630 ;
        RECT 86.935 104.780 87.165 109.930 ;
        RECT 89.225 104.780 89.455 111.430 ;
        RECT 90.565 106.130 90.795 112.780 ;
        RECT 90.330 105.430 91.030 106.130 ;
        RECT 90.565 104.780 90.795 105.430 ;
        RECT 72.805 103.885 77.615 104.780 ;
        RECT 92.855 104.575 93.085 112.780 ;
        RECT 95.145 106.130 95.375 112.780 ;
        RECT 96.485 112.130 96.715 112.780 ;
        RECT 96.250 111.430 96.950 112.130 ;
        RECT 94.910 105.430 95.610 106.130 ;
        RECT 95.145 104.780 95.375 105.430 ;
        RECT 96.485 104.780 96.715 111.430 ;
        RECT 98.775 110.630 99.005 112.780 ;
        RECT 101.065 112.130 101.295 112.780 ;
        RECT 100.830 111.430 101.530 112.130 ;
        RECT 98.540 109.930 99.240 110.630 ;
        RECT 98.775 104.780 99.005 109.930 ;
        RECT 101.065 104.780 101.295 111.430 ;
        RECT 102.405 107.630 102.635 112.780 ;
        RECT 104.695 109.130 104.925 112.780 ;
        RECT 104.460 108.430 105.160 109.130 ;
        RECT 102.170 106.930 102.870 107.630 ;
        RECT 102.405 104.780 102.635 106.930 ;
        RECT 104.695 104.780 104.925 108.430 ;
        RECT 106.985 107.630 107.215 112.780 ;
        RECT 106.750 106.930 107.450 107.630 ;
        RECT 106.985 104.780 107.215 106.930 ;
        RECT 108.325 104.780 108.555 112.780 ;
        RECT 110.615 104.780 110.845 112.780 ;
        RECT 112.905 104.780 113.135 112.780 ;
        RECT 79.005 104.275 80.965 104.575 ;
        RECT 81.295 104.275 83.255 104.575 ;
        RECT 84.925 104.275 86.885 104.575 ;
        RECT 87.215 104.275 89.175 104.575 ;
        RECT 90.845 104.275 95.095 104.575 ;
        RECT 96.765 104.275 98.725 104.575 ;
        RECT 99.055 104.275 101.015 104.575 ;
        RECT 102.685 104.275 104.645 104.575 ;
        RECT 104.975 104.275 106.935 104.575 ;
        RECT 108.325 103.885 113.135 104.780 ;
        RECT 113.575 103.885 114.165 123.695 ;
        RECT 128.935 123.505 135.120 124.285 ;
        RECT 138.080 128.380 145.960 128.970 ;
        RECT 138.080 124.680 138.670 128.380 ;
        RECT 139.205 127.290 139.435 127.530 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 139.205 125.530 139.435 125.690 ;
        RECT 140.495 125.530 140.725 128.380 ;
        RECT 143.725 127.920 144.425 127.990 ;
        RECT 143.595 127.690 144.555 127.920 ;
        RECT 141.785 127.290 142.015 127.530 ;
        RECT 141.700 125.690 142.100 127.290 ;
        RECT 143.315 126.865 143.545 127.530 ;
        RECT 143.280 126.165 143.580 126.865 ;
        RECT 141.785 125.530 142.015 125.690 ;
        RECT 143.315 125.370 143.545 126.165 ;
        RECT 139.390 125.140 143.545 125.370 ;
        RECT 144.605 124.680 144.835 127.530 ;
        RECT 145.370 124.680 145.960 128.380 ;
        RECT 138.080 124.090 145.960 124.680 ;
        RECT 71.775 102.705 114.165 103.885 ;
        RECT 115.905 122.915 135.120 123.505 ;
        RECT 115.905 122.475 116.495 122.915 ;
        RECT 115.905 122.245 118.390 122.475 ;
        RECT 115.905 114.185 117.185 122.245 ;
        RECT 118.595 114.235 118.825 122.195 ;
        RECT 119.975 118.645 120.205 122.195 ;
        RECT 120.410 122.010 121.410 122.710 ;
        RECT 121.615 118.645 121.845 122.195 ;
        RECT 119.975 117.075 121.845 118.645 ;
        RECT 115.905 113.955 118.390 114.185 ;
        RECT 115.905 112.845 116.495 113.955 ;
        RECT 115.905 112.615 118.390 112.845 ;
        RECT 115.905 104.555 117.185 112.615 ;
        RECT 118.595 104.605 118.825 112.565 ;
        RECT 119.975 109.685 120.205 117.075 ;
        RECT 121.615 114.235 121.845 117.075 ;
        RECT 122.995 118.645 123.225 122.195 ;
        RECT 123.430 122.010 124.430 122.710 ;
        RECT 128.345 122.475 135.120 122.915 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 126.450 122.245 135.120 122.475 ;
        RECT 124.635 118.645 124.865 122.195 ;
        RECT 122.995 117.075 124.865 118.645 ;
        RECT 122.995 114.235 123.225 117.075 ;
        RECT 120.410 112.615 121.410 114.185 ;
        RECT 123.430 112.615 124.430 114.185 ;
        RECT 121.615 109.685 121.845 112.565 ;
        RECT 119.975 108.115 121.845 109.685 ;
        RECT 119.975 104.605 120.205 108.115 ;
        RECT 115.905 104.325 118.390 104.555 ;
        RECT 115.905 103.885 116.495 104.325 ;
        RECT 120.410 104.090 121.410 104.790 ;
        RECT 121.615 104.605 121.845 108.115 ;
        RECT 122.995 109.685 123.225 112.565 ;
        RECT 124.635 109.685 124.865 117.075 ;
        RECT 126.015 114.235 126.245 122.195 ;
        RECT 127.655 114.185 135.120 122.245 ;
        RECT 126.450 113.955 135.120 114.185 ;
        RECT 128.345 112.845 135.120 113.955 ;
        RECT 126.450 112.615 135.120 112.845 ;
        RECT 122.995 108.115 124.865 109.685 ;
        RECT 122.995 104.605 123.225 108.115 ;
        RECT 123.430 104.090 124.430 104.790 ;
        RECT 124.635 104.605 124.865 108.115 ;
        RECT 126.015 104.605 126.245 112.565 ;
        RECT 127.655 107.765 135.120 112.615 ;
        RECT 136.295 108.925 142.995 109.515 ;
        RECT 127.655 104.835 138.400 107.765 ;
        RECT 127.655 104.555 135.710 104.835 ;
        RECT 126.450 104.325 135.710 104.555 ;
        RECT 128.345 103.885 135.710 104.325 ;
        RECT 115.905 102.705 135.710 103.885 ;
        RECT 8.665 102.115 135.710 102.705 ;
        RECT 136.295 102.495 138.400 104.255 ;
        RECT 8.665 44.835 10.615 102.115 ;
        RECT 4.100 42.225 10.615 44.835 ;
        RECT 11.055 101.425 29.605 102.115 ;
        RECT 11.055 93.015 11.285 101.425 ;
        RECT 13.345 93.015 13.575 101.425 ;
        RECT 15.635 93.015 15.865 101.425 ;
        RECT 17.925 93.015 18.155 101.425 ;
        RECT 20.215 93.015 20.445 101.425 ;
        RECT 22.505 93.015 22.735 101.425 ;
        RECT 24.795 93.015 25.025 101.425 ;
        RECT 27.085 93.015 27.315 101.425 ;
        RECT 29.375 93.015 29.605 101.425 ;
        RECT 30.715 101.425 49.265 102.115 ;
        RECT 30.715 93.220 30.945 101.425 ;
        RECT 33.005 93.220 33.235 101.425 ;
        RECT 35.295 93.220 35.525 101.425 ;
        RECT 37.585 93.220 37.815 101.425 ;
        RECT 39.875 93.220 40.105 101.425 ;
        RECT 42.165 93.220 42.395 101.425 ;
        RECT 44.455 93.220 44.685 101.425 ;
        RECT 46.745 93.220 46.975 101.425 ;
        RECT 49.035 93.220 49.265 101.425 ;
        RECT 50.375 101.425 68.925 102.115 ;
        RECT 50.375 93.220 50.605 101.425 ;
        RECT 52.665 93.220 52.895 101.425 ;
        RECT 54.955 93.220 55.185 101.425 ;
        RECT 57.245 93.220 57.475 101.425 ;
        RECT 59.535 93.220 59.765 101.425 ;
        RECT 61.825 93.220 62.055 101.425 ;
        RECT 64.115 93.220 64.345 101.425 ;
        RECT 66.405 93.220 66.635 101.425 ;
        RECT 68.695 93.220 68.925 101.425 ;
        RECT 70.035 101.425 88.585 102.115 ;
        RECT 70.035 93.220 70.265 101.425 ;
        RECT 72.325 93.220 72.555 101.425 ;
        RECT 74.615 93.220 74.845 101.425 ;
        RECT 76.905 93.220 77.135 101.425 ;
        RECT 79.195 93.220 79.425 101.425 ;
        RECT 81.485 93.220 81.715 101.425 ;
        RECT 83.775 93.220 84.005 101.425 ;
        RECT 86.065 93.220 86.295 101.425 ;
        RECT 88.355 93.220 88.585 101.425 ;
        RECT 89.695 101.425 108.245 102.115 ;
        RECT 89.695 93.220 89.925 101.425 ;
        RECT 91.985 93.220 92.215 101.425 ;
        RECT 94.275 93.220 94.505 101.425 ;
        RECT 96.565 93.220 96.795 101.425 ;
        RECT 98.855 93.220 99.085 101.425 ;
        RECT 101.145 93.220 101.375 101.425 ;
        RECT 103.435 93.220 103.665 101.425 ;
        RECT 105.725 93.220 105.955 101.425 ;
        RECT 108.015 93.220 108.245 101.425 ;
        RECT 109.355 101.425 127.905 102.115 ;
        RECT 109.355 93.015 109.585 101.425 ;
        RECT 111.645 93.015 111.875 101.425 ;
        RECT 113.935 93.015 114.165 101.425 ;
        RECT 116.225 93.015 116.455 101.425 ;
        RECT 118.515 93.015 118.745 101.425 ;
        RECT 120.805 93.015 121.035 101.425 ;
        RECT 123.095 93.015 123.325 101.425 ;
        RECT 125.385 93.015 125.615 101.425 ;
        RECT 127.675 93.015 127.905 101.425 ;
        RECT 11.055 91.405 29.605 93.015 ;
        RECT 30.995 92.785 32.955 93.015 ;
        RECT 33.285 92.785 35.245 93.015 ;
        RECT 35.575 92.785 37.535 93.015 ;
        RECT 37.865 92.785 39.825 93.015 ;
        RECT 40.155 92.785 42.115 93.015 ;
        RECT 42.445 92.785 44.405 93.015 ;
        RECT 44.735 92.785 46.695 93.015 ;
        RECT 47.025 92.785 48.985 93.015 ;
        RECT 50.655 92.785 52.615 93.015 ;
        RECT 52.945 92.785 54.905 93.015 ;
        RECT 55.235 92.785 57.195 93.015 ;
        RECT 57.525 92.785 59.485 93.015 ;
        RECT 59.815 92.785 61.775 93.015 ;
        RECT 62.105 92.785 64.065 93.015 ;
        RECT 64.395 92.785 66.355 93.015 ;
        RECT 66.685 92.785 68.645 93.015 ;
        RECT 70.315 92.785 72.275 93.015 ;
        RECT 72.605 92.785 74.565 93.015 ;
        RECT 74.895 92.785 76.855 93.015 ;
        RECT 77.185 92.785 79.145 93.015 ;
        RECT 79.475 92.785 81.435 93.015 ;
        RECT 81.765 92.785 83.725 93.015 ;
        RECT 84.055 92.785 86.015 93.015 ;
        RECT 86.345 92.785 88.305 93.015 ;
        RECT 89.975 92.785 91.935 93.015 ;
        RECT 92.265 92.785 94.225 93.015 ;
        RECT 94.555 92.785 96.515 93.015 ;
        RECT 96.845 92.785 98.805 93.015 ;
        RECT 99.135 92.785 101.095 93.015 ;
        RECT 101.425 92.785 103.385 93.015 ;
        RECT 103.715 92.785 105.675 93.015 ;
        RECT 106.005 92.785 107.965 93.015 ;
        RECT 30.995 91.405 32.955 91.635 ;
        RECT 11.055 82.995 11.285 91.405 ;
        RECT 13.345 82.995 13.575 91.405 ;
        RECT 15.635 82.995 15.865 91.405 ;
        RECT 17.925 82.995 18.155 91.405 ;
        RECT 20.215 82.995 20.445 91.405 ;
        RECT 22.505 82.995 22.735 91.405 ;
        RECT 24.795 82.995 25.025 91.405 ;
        RECT 27.085 82.995 27.315 91.405 ;
        RECT 29.375 82.995 29.605 91.405 ;
        RECT 33.285 91.345 35.245 91.875 ;
        RECT 35.575 91.345 37.535 91.875 ;
        RECT 37.865 91.405 39.825 91.635 ;
        RECT 40.155 91.405 42.115 91.635 ;
        RECT 42.445 91.345 44.405 91.875 ;
        RECT 44.735 91.345 46.695 91.875 ;
        RECT 47.025 91.405 48.985 91.635 ;
        RECT 50.655 91.345 52.615 91.875 ;
        RECT 52.945 91.405 54.905 91.635 ;
        RECT 55.235 91.405 57.195 91.635 ;
        RECT 57.525 91.345 59.485 91.875 ;
        RECT 59.815 91.345 61.775 91.875 ;
        RECT 62.105 91.405 64.065 91.635 ;
        RECT 64.395 91.405 66.355 91.635 ;
        RECT 66.685 91.345 68.645 91.875 ;
        RECT 70.315 91.345 72.275 91.875 ;
        RECT 72.605 91.405 74.565 91.635 ;
        RECT 74.895 91.405 76.855 91.635 ;
        RECT 77.185 91.345 79.145 91.875 ;
        RECT 79.475 91.345 81.435 91.875 ;
        RECT 81.765 91.405 83.725 91.635 ;
        RECT 84.055 91.405 86.015 91.635 ;
        RECT 86.345 91.345 88.305 91.875 ;
        RECT 89.975 91.405 91.935 91.635 ;
        RECT 92.265 91.345 94.225 91.875 ;
        RECT 94.555 91.345 96.515 91.875 ;
        RECT 96.845 91.405 98.805 91.635 ;
        RECT 99.135 91.405 101.095 91.635 ;
        RECT 101.425 91.345 103.385 91.875 ;
        RECT 103.715 91.345 105.675 91.875 ;
        RECT 106.005 91.405 107.965 91.635 ;
        RECT 109.355 91.405 127.905 93.015 ;
        RECT 30.715 84.590 30.945 91.200 ;
        RECT 33.005 88.540 33.235 91.200 ;
        RECT 35.295 91.090 35.525 91.200 ;
        RECT 35.260 89.690 35.560 91.090 ;
        RECT 32.970 85.740 33.270 88.540 ;
        RECT 30.680 83.190 30.980 84.590 ;
        RECT 33.005 83.200 33.235 85.740 ;
        RECT 35.295 83.200 35.525 89.690 ;
        RECT 37.585 88.540 37.815 91.200 ;
        RECT 37.550 85.740 37.850 88.540 ;
        RECT 37.585 83.200 37.815 85.740 ;
        RECT 39.875 84.590 40.105 91.200 ;
        RECT 42.165 88.540 42.395 91.200 ;
        RECT 44.455 91.090 44.685 91.200 ;
        RECT 44.420 89.690 44.720 91.090 ;
        RECT 42.130 85.740 42.430 88.540 ;
        RECT 39.840 83.190 40.140 84.590 ;
        RECT 42.165 83.200 42.395 85.740 ;
        RECT 44.455 83.200 44.685 89.690 ;
        RECT 46.745 88.540 46.975 91.200 ;
        RECT 46.710 85.740 47.010 88.540 ;
        RECT 46.745 83.200 46.975 85.740 ;
        RECT 49.035 84.590 49.265 91.200 ;
        RECT 50.375 91.090 50.605 91.200 ;
        RECT 50.340 89.690 50.640 91.090 ;
        RECT 49.000 83.190 49.300 84.590 ;
        RECT 50.375 83.200 50.605 89.690 ;
        RECT 52.665 88.540 52.895 91.200 ;
        RECT 52.630 85.740 52.930 88.540 ;
        RECT 52.665 83.200 52.895 85.740 ;
        RECT 54.955 84.590 55.185 91.200 ;
        RECT 57.245 88.540 57.475 91.200 ;
        RECT 59.535 91.090 59.765 91.200 ;
        RECT 59.500 89.690 59.800 91.090 ;
        RECT 57.210 85.740 57.510 88.540 ;
        RECT 54.920 83.190 55.220 84.590 ;
        RECT 57.245 83.200 57.475 85.740 ;
        RECT 59.535 83.200 59.765 89.690 ;
        RECT 61.825 88.540 62.055 91.200 ;
        RECT 61.790 85.740 62.090 88.540 ;
        RECT 61.825 83.200 62.055 85.740 ;
        RECT 64.115 84.590 64.345 91.200 ;
        RECT 66.405 88.540 66.635 91.200 ;
        RECT 68.695 91.090 68.925 91.200 ;
        RECT 70.035 91.090 70.265 91.200 ;
        RECT 68.660 89.690 68.960 91.090 ;
        RECT 70.000 89.690 70.300 91.090 ;
        RECT 66.370 85.740 66.670 88.540 ;
        RECT 64.080 83.190 64.380 84.590 ;
        RECT 66.405 83.200 66.635 85.740 ;
        RECT 68.695 83.200 68.925 89.690 ;
        RECT 70.035 83.200 70.265 89.690 ;
        RECT 72.325 88.540 72.555 91.200 ;
        RECT 72.290 85.740 72.590 88.540 ;
        RECT 72.325 83.200 72.555 85.740 ;
        RECT 74.615 84.590 74.845 91.200 ;
        RECT 76.905 88.540 77.135 91.200 ;
        RECT 79.195 91.090 79.425 91.200 ;
        RECT 79.160 89.690 79.460 91.090 ;
        RECT 76.870 85.740 77.170 88.540 ;
        RECT 74.580 83.190 74.880 84.590 ;
        RECT 76.905 83.200 77.135 85.740 ;
        RECT 79.195 83.200 79.425 89.690 ;
        RECT 81.485 88.540 81.715 91.200 ;
        RECT 81.450 85.740 81.750 88.540 ;
        RECT 81.485 83.200 81.715 85.740 ;
        RECT 83.775 84.590 84.005 91.200 ;
        RECT 86.065 88.540 86.295 91.200 ;
        RECT 88.355 91.090 88.585 91.200 ;
        RECT 88.320 89.690 88.620 91.090 ;
        RECT 86.030 85.740 86.330 88.540 ;
        RECT 83.740 83.190 84.040 84.590 ;
        RECT 86.065 83.200 86.295 85.740 ;
        RECT 88.355 83.200 88.585 89.690 ;
        RECT 89.695 84.590 89.925 91.200 ;
        RECT 91.985 88.540 92.215 91.200 ;
        RECT 94.275 91.090 94.505 91.200 ;
        RECT 94.240 89.690 94.540 91.090 ;
        RECT 91.950 85.740 92.250 88.540 ;
        RECT 89.660 83.190 89.960 84.590 ;
        RECT 91.985 83.200 92.215 85.740 ;
        RECT 94.275 83.200 94.505 89.690 ;
        RECT 96.565 88.540 96.795 91.200 ;
        RECT 96.530 85.740 96.830 88.540 ;
        RECT 96.565 83.200 96.795 85.740 ;
        RECT 98.855 84.590 99.085 91.200 ;
        RECT 101.145 88.540 101.375 91.200 ;
        RECT 103.435 91.090 103.665 91.200 ;
        RECT 103.400 89.690 103.700 91.090 ;
        RECT 101.110 85.740 101.410 88.540 ;
        RECT 98.820 83.190 99.120 84.590 ;
        RECT 101.145 83.200 101.375 85.740 ;
        RECT 103.435 83.200 103.665 89.690 ;
        RECT 105.725 88.540 105.955 91.200 ;
        RECT 105.690 85.740 105.990 88.540 ;
        RECT 105.725 83.200 105.955 85.740 ;
        RECT 108.015 84.590 108.245 91.200 ;
        RECT 107.980 83.190 108.280 84.590 ;
        RECT 109.355 82.995 109.585 91.405 ;
        RECT 111.645 82.995 111.875 91.405 ;
        RECT 113.935 82.995 114.165 91.405 ;
        RECT 116.225 82.995 116.455 91.405 ;
        RECT 118.515 82.995 118.745 91.405 ;
        RECT 120.805 82.995 121.035 91.405 ;
        RECT 123.095 82.995 123.325 91.405 ;
        RECT 125.385 82.995 125.615 91.405 ;
        RECT 127.675 82.995 127.905 91.405 ;
        RECT 11.055 81.385 29.605 82.995 ;
        RECT 30.995 82.405 32.955 82.995 ;
        RECT 33.285 82.765 35.245 82.995 ;
        RECT 35.575 82.765 37.535 82.995 ;
        RECT 37.865 82.405 39.825 82.995 ;
        RECT 40.155 82.405 42.115 82.995 ;
        RECT 42.445 82.765 44.405 82.995 ;
        RECT 44.735 82.765 46.695 82.995 ;
        RECT 47.025 82.405 48.985 82.995 ;
        RECT 50.655 82.765 52.615 82.995 ;
        RECT 52.945 82.405 54.905 82.995 ;
        RECT 55.235 82.405 57.195 82.995 ;
        RECT 57.525 82.765 59.485 82.995 ;
        RECT 59.815 82.765 61.775 82.995 ;
        RECT 62.105 82.405 64.065 82.995 ;
        RECT 64.395 82.405 66.355 82.995 ;
        RECT 66.685 82.765 68.645 82.995 ;
        RECT 70.315 82.765 72.275 82.995 ;
        RECT 72.605 82.405 74.565 82.995 ;
        RECT 74.895 82.405 76.855 82.995 ;
        RECT 77.185 82.765 79.145 82.995 ;
        RECT 79.475 82.765 81.435 82.995 ;
        RECT 81.765 82.405 83.725 82.995 ;
        RECT 84.055 82.405 86.015 82.995 ;
        RECT 86.345 82.765 88.305 82.995 ;
        RECT 89.975 82.405 91.935 82.995 ;
        RECT 92.265 82.765 94.225 82.995 ;
        RECT 94.555 82.765 96.515 82.995 ;
        RECT 96.845 82.405 98.805 82.995 ;
        RECT 99.135 82.405 101.095 82.995 ;
        RECT 101.425 82.765 103.385 82.995 ;
        RECT 103.715 82.765 105.675 82.995 ;
        RECT 106.005 82.405 107.965 82.995 ;
        RECT 30.995 81.385 32.955 81.615 ;
        RECT 11.055 72.975 11.285 81.385 ;
        RECT 13.345 72.975 13.575 81.385 ;
        RECT 15.635 72.975 15.865 81.385 ;
        RECT 17.925 72.975 18.155 81.385 ;
        RECT 20.215 72.975 20.445 81.385 ;
        RECT 22.505 72.975 22.735 81.385 ;
        RECT 24.795 72.975 25.025 81.385 ;
        RECT 27.085 72.975 27.315 81.385 ;
        RECT 29.375 72.975 29.605 81.385 ;
        RECT 33.285 81.325 35.245 81.855 ;
        RECT 35.575 81.325 37.535 81.855 ;
        RECT 37.865 81.385 39.825 81.615 ;
        RECT 40.155 81.385 42.115 81.615 ;
        RECT 42.445 81.325 44.405 81.855 ;
        RECT 44.735 81.325 46.695 81.855 ;
        RECT 47.025 81.385 48.985 81.615 ;
        RECT 50.655 81.325 52.615 81.855 ;
        RECT 52.945 81.385 54.905 81.615 ;
        RECT 55.235 81.385 57.195 81.615 ;
        RECT 57.525 81.325 59.485 81.855 ;
        RECT 59.815 81.325 61.775 81.855 ;
        RECT 62.105 81.385 64.065 81.615 ;
        RECT 64.395 81.385 66.355 81.615 ;
        RECT 66.685 81.325 68.645 81.855 ;
        RECT 70.315 81.325 72.275 81.855 ;
        RECT 72.605 81.385 74.565 81.615 ;
        RECT 74.895 81.385 76.855 81.615 ;
        RECT 77.185 81.325 79.145 81.855 ;
        RECT 79.475 81.325 81.435 81.855 ;
        RECT 81.765 81.385 83.725 81.615 ;
        RECT 84.055 81.385 86.015 81.615 ;
        RECT 86.345 81.325 88.305 81.855 ;
        RECT 89.975 81.385 91.935 81.615 ;
        RECT 92.265 81.325 94.225 81.855 ;
        RECT 94.555 81.325 96.515 81.855 ;
        RECT 96.845 81.385 98.805 81.615 ;
        RECT 99.135 81.385 101.095 81.615 ;
        RECT 101.425 81.325 103.385 81.855 ;
        RECT 103.715 81.325 105.675 81.855 ;
        RECT 106.005 81.385 107.965 81.615 ;
        RECT 109.355 81.385 127.905 82.995 ;
        RECT 30.715 81.070 30.945 81.180 ;
        RECT 30.680 79.670 30.980 81.070 ;
        RECT 30.715 73.180 30.945 79.670 ;
        RECT 33.005 78.520 33.235 81.180 ;
        RECT 32.970 75.720 33.270 78.520 ;
        RECT 33.005 73.180 33.235 75.720 ;
        RECT 35.295 74.570 35.525 81.180 ;
        RECT 37.585 78.520 37.815 81.180 ;
        RECT 39.875 81.070 40.105 81.180 ;
        RECT 39.840 79.670 40.140 81.070 ;
        RECT 37.550 75.720 37.850 78.520 ;
        RECT 35.260 73.170 35.560 74.570 ;
        RECT 37.585 73.180 37.815 75.720 ;
        RECT 39.875 73.180 40.105 79.670 ;
        RECT 42.165 78.520 42.395 81.180 ;
        RECT 42.130 75.720 42.430 78.520 ;
        RECT 42.165 73.180 42.395 75.720 ;
        RECT 44.455 74.570 44.685 81.180 ;
        RECT 46.745 78.520 46.975 81.180 ;
        RECT 49.035 81.070 49.265 81.180 ;
        RECT 49.000 79.670 49.300 81.070 ;
        RECT 46.710 75.720 47.010 78.520 ;
        RECT 44.420 73.170 44.720 74.570 ;
        RECT 46.745 73.180 46.975 75.720 ;
        RECT 49.035 73.180 49.265 79.670 ;
        RECT 50.375 74.570 50.605 81.180 ;
        RECT 52.665 78.520 52.895 81.180 ;
        RECT 54.955 81.070 55.185 81.180 ;
        RECT 54.920 79.670 55.220 81.070 ;
        RECT 52.630 75.720 52.930 78.520 ;
        RECT 50.340 73.170 50.640 74.570 ;
        RECT 52.665 73.180 52.895 75.720 ;
        RECT 54.955 73.180 55.185 79.670 ;
        RECT 57.245 78.520 57.475 81.180 ;
        RECT 57.210 75.720 57.510 78.520 ;
        RECT 57.245 73.180 57.475 75.720 ;
        RECT 59.535 74.570 59.765 81.180 ;
        RECT 61.825 78.520 62.055 81.180 ;
        RECT 64.115 81.070 64.345 81.180 ;
        RECT 64.080 79.670 64.380 81.070 ;
        RECT 61.790 75.720 62.090 78.520 ;
        RECT 59.500 73.170 59.800 74.570 ;
        RECT 61.825 73.180 62.055 75.720 ;
        RECT 64.115 73.180 64.345 79.670 ;
        RECT 66.405 78.520 66.635 81.180 ;
        RECT 66.370 75.720 66.670 78.520 ;
        RECT 66.405 73.180 66.635 75.720 ;
        RECT 68.695 74.570 68.925 81.180 ;
        RECT 70.035 74.570 70.265 81.180 ;
        RECT 72.325 78.520 72.555 81.180 ;
        RECT 74.615 81.070 74.845 81.180 ;
        RECT 74.580 79.670 74.880 81.070 ;
        RECT 72.290 75.720 72.590 78.520 ;
        RECT 68.660 73.170 68.960 74.570 ;
        RECT 70.000 73.170 70.300 74.570 ;
        RECT 72.325 73.180 72.555 75.720 ;
        RECT 74.615 73.180 74.845 79.670 ;
        RECT 76.905 78.520 77.135 81.180 ;
        RECT 76.870 75.720 77.170 78.520 ;
        RECT 76.905 73.180 77.135 75.720 ;
        RECT 79.195 74.570 79.425 81.180 ;
        RECT 81.485 78.520 81.715 81.180 ;
        RECT 83.775 81.070 84.005 81.180 ;
        RECT 83.740 79.670 84.040 81.070 ;
        RECT 81.450 75.720 81.750 78.520 ;
        RECT 79.160 73.170 79.460 74.570 ;
        RECT 81.485 73.180 81.715 75.720 ;
        RECT 83.775 73.180 84.005 79.670 ;
        RECT 86.065 78.520 86.295 81.180 ;
        RECT 86.030 75.720 86.330 78.520 ;
        RECT 86.065 73.180 86.295 75.720 ;
        RECT 88.355 74.570 88.585 81.180 ;
        RECT 89.695 81.070 89.925 81.180 ;
        RECT 89.660 79.670 89.960 81.070 ;
        RECT 88.320 73.170 88.620 74.570 ;
        RECT 89.695 73.180 89.925 79.670 ;
        RECT 91.985 78.520 92.215 81.180 ;
        RECT 91.950 75.720 92.250 78.520 ;
        RECT 91.985 73.180 92.215 75.720 ;
        RECT 94.275 74.570 94.505 81.180 ;
        RECT 96.565 78.520 96.795 81.180 ;
        RECT 98.855 81.070 99.085 81.180 ;
        RECT 98.820 79.670 99.120 81.070 ;
        RECT 96.530 75.720 96.830 78.520 ;
        RECT 94.240 73.170 94.540 74.570 ;
        RECT 96.565 73.180 96.795 75.720 ;
        RECT 98.855 73.180 99.085 79.670 ;
        RECT 101.145 78.520 101.375 81.180 ;
        RECT 101.110 75.720 101.410 78.520 ;
        RECT 101.145 73.180 101.375 75.720 ;
        RECT 103.435 74.570 103.665 81.180 ;
        RECT 105.725 78.520 105.955 81.180 ;
        RECT 108.015 81.070 108.245 81.180 ;
        RECT 107.980 79.670 108.280 81.070 ;
        RECT 105.690 75.720 105.990 78.520 ;
        RECT 103.400 73.170 103.700 74.570 ;
        RECT 105.725 73.180 105.955 75.720 ;
        RECT 108.015 73.180 108.245 79.670 ;
        RECT 109.355 72.975 109.585 81.385 ;
        RECT 111.645 72.975 111.875 81.385 ;
        RECT 113.935 72.975 114.165 81.385 ;
        RECT 116.225 72.975 116.455 81.385 ;
        RECT 118.515 72.975 118.745 81.385 ;
        RECT 120.805 72.975 121.035 81.385 ;
        RECT 123.095 72.975 123.325 81.385 ;
        RECT 125.385 72.975 125.615 81.385 ;
        RECT 127.675 72.975 127.905 81.385 ;
        RECT 11.055 71.365 29.605 72.975 ;
        RECT 30.995 72.385 32.955 72.975 ;
        RECT 33.285 72.745 35.245 72.975 ;
        RECT 35.575 72.745 37.535 72.975 ;
        RECT 37.865 72.385 39.825 72.975 ;
        RECT 40.155 72.385 42.115 72.975 ;
        RECT 42.445 72.745 44.405 72.975 ;
        RECT 44.735 72.745 46.695 72.975 ;
        RECT 47.025 72.385 48.985 72.975 ;
        RECT 50.655 72.745 52.615 72.975 ;
        RECT 52.945 72.385 54.905 72.975 ;
        RECT 55.235 72.385 57.195 72.975 ;
        RECT 57.525 72.745 59.485 72.975 ;
        RECT 59.815 72.745 61.775 72.975 ;
        RECT 62.105 72.385 64.065 72.975 ;
        RECT 64.395 72.385 66.355 72.975 ;
        RECT 66.685 72.745 68.645 72.975 ;
        RECT 70.315 72.745 72.275 72.975 ;
        RECT 72.605 72.385 74.565 72.975 ;
        RECT 74.895 72.385 76.855 72.975 ;
        RECT 77.185 72.745 79.145 72.975 ;
        RECT 79.475 72.745 81.435 72.975 ;
        RECT 81.765 72.385 83.725 72.975 ;
        RECT 84.055 72.385 86.015 72.975 ;
        RECT 86.345 72.745 88.305 72.975 ;
        RECT 89.975 72.385 91.935 72.975 ;
        RECT 92.265 72.745 94.225 72.975 ;
        RECT 94.555 72.745 96.515 72.975 ;
        RECT 96.845 72.385 98.805 72.975 ;
        RECT 99.135 72.385 101.095 72.975 ;
        RECT 101.425 72.745 103.385 72.975 ;
        RECT 103.715 72.745 105.675 72.975 ;
        RECT 106.005 72.385 107.965 72.975 ;
        RECT 11.055 62.955 11.285 71.365 ;
        RECT 13.345 62.955 13.575 71.365 ;
        RECT 15.635 62.955 15.865 71.365 ;
        RECT 17.925 62.955 18.155 71.365 ;
        RECT 20.215 62.955 20.445 71.365 ;
        RECT 22.505 62.955 22.735 71.365 ;
        RECT 24.795 62.955 25.025 71.365 ;
        RECT 27.085 62.955 27.315 71.365 ;
        RECT 29.375 62.955 29.605 71.365 ;
        RECT 30.995 71.305 32.955 71.835 ;
        RECT 33.285 71.365 35.245 71.595 ;
        RECT 35.575 71.365 37.535 71.595 ;
        RECT 37.865 71.305 39.825 71.835 ;
        RECT 40.155 71.305 42.115 71.835 ;
        RECT 42.445 71.365 44.405 71.595 ;
        RECT 44.735 71.365 46.695 71.595 ;
        RECT 47.025 71.305 48.985 71.835 ;
        RECT 50.655 71.365 52.615 71.595 ;
        RECT 52.945 71.305 54.905 71.835 ;
        RECT 55.235 71.305 57.195 71.835 ;
        RECT 57.525 71.365 59.485 71.595 ;
        RECT 59.815 71.365 61.775 71.595 ;
        RECT 62.105 71.305 64.065 71.835 ;
        RECT 64.395 71.305 66.355 71.835 ;
        RECT 66.685 71.365 68.645 71.595 ;
        RECT 70.315 71.365 72.275 71.595 ;
        RECT 72.605 71.305 74.565 71.835 ;
        RECT 74.895 71.305 76.855 71.835 ;
        RECT 77.185 71.365 79.145 71.595 ;
        RECT 79.475 71.365 81.435 71.595 ;
        RECT 81.765 71.305 83.725 71.835 ;
        RECT 84.055 71.305 86.015 71.835 ;
        RECT 86.345 71.365 88.305 71.595 ;
        RECT 89.975 71.305 91.935 71.835 ;
        RECT 92.265 71.365 94.225 71.595 ;
        RECT 94.555 71.365 96.515 71.595 ;
        RECT 96.845 71.305 98.805 71.835 ;
        RECT 99.135 71.305 101.095 71.835 ;
        RECT 101.425 71.365 103.385 71.595 ;
        RECT 103.715 71.365 105.675 71.595 ;
        RECT 106.005 71.305 107.965 71.835 ;
        RECT 109.355 71.365 127.905 72.975 ;
        RECT 30.715 71.050 30.945 71.160 ;
        RECT 30.680 69.650 30.980 71.050 ;
        RECT 30.715 63.160 30.945 69.650 ;
        RECT 33.005 68.500 33.235 71.160 ;
        RECT 32.970 65.700 33.270 68.500 ;
        RECT 33.005 63.160 33.235 65.700 ;
        RECT 35.295 64.550 35.525 71.160 ;
        RECT 37.585 68.500 37.815 71.160 ;
        RECT 39.875 71.050 40.105 71.160 ;
        RECT 39.840 69.650 40.140 71.050 ;
        RECT 37.550 65.700 37.850 68.500 ;
        RECT 35.260 63.150 35.560 64.550 ;
        RECT 37.585 63.160 37.815 65.700 ;
        RECT 39.875 63.160 40.105 69.650 ;
        RECT 42.165 68.500 42.395 71.160 ;
        RECT 42.130 65.700 42.430 68.500 ;
        RECT 42.165 63.160 42.395 65.700 ;
        RECT 44.455 64.550 44.685 71.160 ;
        RECT 46.745 68.500 46.975 71.160 ;
        RECT 49.035 71.050 49.265 71.160 ;
        RECT 49.000 69.650 49.300 71.050 ;
        RECT 46.710 65.700 47.010 68.500 ;
        RECT 44.420 63.150 44.720 64.550 ;
        RECT 46.745 63.160 46.975 65.700 ;
        RECT 49.035 63.160 49.265 69.650 ;
        RECT 50.375 64.550 50.605 71.160 ;
        RECT 52.665 68.500 52.895 71.160 ;
        RECT 54.955 71.050 55.185 71.160 ;
        RECT 54.920 69.650 55.220 71.050 ;
        RECT 52.630 65.700 52.930 68.500 ;
        RECT 50.340 63.150 50.640 64.550 ;
        RECT 52.665 63.160 52.895 65.700 ;
        RECT 54.955 63.160 55.185 69.650 ;
        RECT 57.245 68.500 57.475 71.160 ;
        RECT 57.210 65.700 57.510 68.500 ;
        RECT 57.245 63.160 57.475 65.700 ;
        RECT 59.535 64.550 59.765 71.160 ;
        RECT 61.825 68.500 62.055 71.160 ;
        RECT 64.115 71.050 64.345 71.160 ;
        RECT 64.080 69.650 64.380 71.050 ;
        RECT 61.790 65.700 62.090 68.500 ;
        RECT 59.500 63.150 59.800 64.550 ;
        RECT 61.825 63.160 62.055 65.700 ;
        RECT 64.115 63.160 64.345 69.650 ;
        RECT 66.405 68.500 66.635 71.160 ;
        RECT 66.370 65.700 66.670 68.500 ;
        RECT 66.405 63.160 66.635 65.700 ;
        RECT 68.695 64.550 68.925 71.160 ;
        RECT 70.035 64.550 70.265 71.160 ;
        RECT 72.325 68.500 72.555 71.160 ;
        RECT 74.615 71.050 74.845 71.160 ;
        RECT 74.580 69.650 74.880 71.050 ;
        RECT 72.290 65.700 72.590 68.500 ;
        RECT 68.660 63.150 68.960 64.550 ;
        RECT 70.000 63.150 70.300 64.550 ;
        RECT 72.325 63.160 72.555 65.700 ;
        RECT 74.615 63.160 74.845 69.650 ;
        RECT 76.905 68.500 77.135 71.160 ;
        RECT 76.870 65.700 77.170 68.500 ;
        RECT 76.905 63.160 77.135 65.700 ;
        RECT 79.195 64.550 79.425 71.160 ;
        RECT 81.485 68.500 81.715 71.160 ;
        RECT 83.775 71.050 84.005 71.160 ;
        RECT 83.740 69.650 84.040 71.050 ;
        RECT 81.450 65.700 81.750 68.500 ;
        RECT 79.160 63.150 79.460 64.550 ;
        RECT 81.485 63.160 81.715 65.700 ;
        RECT 83.775 63.160 84.005 69.650 ;
        RECT 86.065 68.500 86.295 71.160 ;
        RECT 86.030 65.700 86.330 68.500 ;
        RECT 86.065 63.160 86.295 65.700 ;
        RECT 88.355 64.550 88.585 71.160 ;
        RECT 89.695 71.050 89.925 71.160 ;
        RECT 89.660 69.650 89.960 71.050 ;
        RECT 88.320 63.150 88.620 64.550 ;
        RECT 89.695 63.160 89.925 69.650 ;
        RECT 91.985 68.500 92.215 71.160 ;
        RECT 91.950 65.700 92.250 68.500 ;
        RECT 91.985 63.160 92.215 65.700 ;
        RECT 94.275 64.550 94.505 71.160 ;
        RECT 96.565 68.500 96.795 71.160 ;
        RECT 98.855 71.050 99.085 71.160 ;
        RECT 98.820 69.650 99.120 71.050 ;
        RECT 96.530 65.700 96.830 68.500 ;
        RECT 94.240 63.150 94.540 64.550 ;
        RECT 96.565 63.160 96.795 65.700 ;
        RECT 98.855 63.160 99.085 69.650 ;
        RECT 101.145 68.500 101.375 71.160 ;
        RECT 101.110 65.700 101.410 68.500 ;
        RECT 101.145 63.160 101.375 65.700 ;
        RECT 103.435 64.550 103.665 71.160 ;
        RECT 105.725 68.500 105.955 71.160 ;
        RECT 108.015 71.050 108.245 71.160 ;
        RECT 107.980 69.650 108.280 71.050 ;
        RECT 105.690 65.700 105.990 68.500 ;
        RECT 103.400 63.150 103.700 64.550 ;
        RECT 105.725 63.160 105.955 65.700 ;
        RECT 108.015 63.160 108.245 69.650 ;
        RECT 109.355 62.955 109.585 71.365 ;
        RECT 111.645 62.955 111.875 71.365 ;
        RECT 113.935 62.955 114.165 71.365 ;
        RECT 116.225 62.955 116.455 71.365 ;
        RECT 118.515 62.955 118.745 71.365 ;
        RECT 120.805 62.955 121.035 71.365 ;
        RECT 123.095 62.955 123.325 71.365 ;
        RECT 125.385 62.955 125.615 71.365 ;
        RECT 127.675 62.955 127.905 71.365 ;
        RECT 11.055 61.345 29.605 62.955 ;
        RECT 30.995 62.725 32.955 62.955 ;
        RECT 33.285 62.365 35.245 62.955 ;
        RECT 35.575 62.365 37.535 62.955 ;
        RECT 37.865 62.725 39.825 62.955 ;
        RECT 40.155 62.725 42.115 62.955 ;
        RECT 42.445 62.365 44.405 62.955 ;
        RECT 44.735 62.365 46.695 62.955 ;
        RECT 47.025 62.725 48.985 62.955 ;
        RECT 50.655 62.365 52.615 62.955 ;
        RECT 52.945 62.725 54.905 62.955 ;
        RECT 55.235 62.725 57.195 62.955 ;
        RECT 57.525 62.365 59.485 62.955 ;
        RECT 59.815 62.365 61.775 62.955 ;
        RECT 62.105 62.725 64.065 62.955 ;
        RECT 64.395 62.725 66.355 62.955 ;
        RECT 66.685 62.365 68.645 62.955 ;
        RECT 70.315 62.365 72.275 62.955 ;
        RECT 72.605 62.725 74.565 62.955 ;
        RECT 74.895 62.725 76.855 62.955 ;
        RECT 77.185 62.365 79.145 62.955 ;
        RECT 79.475 62.365 81.435 62.955 ;
        RECT 81.765 62.725 83.725 62.955 ;
        RECT 84.055 62.725 86.015 62.955 ;
        RECT 86.345 62.365 88.305 62.955 ;
        RECT 89.975 62.725 91.935 62.955 ;
        RECT 92.265 62.365 94.225 62.955 ;
        RECT 94.555 62.365 96.515 62.955 ;
        RECT 96.845 62.725 98.805 62.955 ;
        RECT 99.135 62.725 101.095 62.955 ;
        RECT 101.425 62.365 103.385 62.955 ;
        RECT 103.715 62.365 105.675 62.955 ;
        RECT 106.005 62.725 107.965 62.955 ;
        RECT 11.055 52.935 11.285 61.345 ;
        RECT 13.345 52.935 13.575 61.345 ;
        RECT 15.635 52.935 15.865 61.345 ;
        RECT 17.925 52.935 18.155 61.345 ;
        RECT 20.215 52.935 20.445 61.345 ;
        RECT 22.505 52.935 22.735 61.345 ;
        RECT 24.795 52.935 25.025 61.345 ;
        RECT 27.085 52.935 27.315 61.345 ;
        RECT 29.375 52.935 29.605 61.345 ;
        RECT 30.995 61.285 32.955 61.815 ;
        RECT 33.285 61.345 35.245 61.575 ;
        RECT 35.575 61.345 37.535 61.575 ;
        RECT 37.865 61.285 39.825 61.815 ;
        RECT 40.155 61.285 42.115 61.815 ;
        RECT 42.445 61.345 44.405 61.575 ;
        RECT 44.735 61.345 46.695 61.575 ;
        RECT 47.025 61.285 48.985 61.815 ;
        RECT 50.655 61.345 52.615 61.575 ;
        RECT 52.945 61.285 54.905 61.815 ;
        RECT 55.235 61.285 57.195 61.815 ;
        RECT 57.525 61.345 59.485 61.575 ;
        RECT 59.815 61.345 61.775 61.575 ;
        RECT 62.105 61.285 64.065 61.815 ;
        RECT 64.395 61.285 66.355 61.815 ;
        RECT 66.685 61.345 68.645 61.575 ;
        RECT 70.315 61.345 72.275 61.575 ;
        RECT 72.605 61.285 74.565 61.815 ;
        RECT 74.895 61.285 76.855 61.815 ;
        RECT 77.185 61.345 79.145 61.575 ;
        RECT 79.475 61.345 81.435 61.575 ;
        RECT 81.765 61.285 83.725 61.815 ;
        RECT 84.055 61.285 86.015 61.815 ;
        RECT 86.345 61.345 88.305 61.575 ;
        RECT 89.975 61.285 91.935 61.815 ;
        RECT 92.265 61.345 94.225 61.575 ;
        RECT 94.555 61.345 96.515 61.575 ;
        RECT 96.845 61.285 98.805 61.815 ;
        RECT 99.135 61.285 101.095 61.815 ;
        RECT 101.425 61.345 103.385 61.575 ;
        RECT 103.715 61.345 105.675 61.575 ;
        RECT 106.005 61.285 107.965 61.815 ;
        RECT 109.355 61.345 127.905 62.955 ;
        RECT 30.715 54.530 30.945 61.140 ;
        RECT 33.005 58.480 33.235 61.140 ;
        RECT 35.295 61.030 35.525 61.140 ;
        RECT 35.260 59.630 35.560 61.030 ;
        RECT 32.970 55.680 33.270 58.480 ;
        RECT 30.680 53.130 30.980 54.530 ;
        RECT 33.005 53.140 33.235 55.680 ;
        RECT 35.295 53.140 35.525 59.630 ;
        RECT 37.585 58.480 37.815 61.140 ;
        RECT 37.550 55.680 37.850 58.480 ;
        RECT 37.585 53.140 37.815 55.680 ;
        RECT 39.875 54.530 40.105 61.140 ;
        RECT 42.165 58.480 42.395 61.140 ;
        RECT 44.455 61.030 44.685 61.140 ;
        RECT 44.420 59.630 44.720 61.030 ;
        RECT 42.130 55.680 42.430 58.480 ;
        RECT 39.840 53.130 40.140 54.530 ;
        RECT 42.165 53.140 42.395 55.680 ;
        RECT 44.455 53.140 44.685 59.630 ;
        RECT 46.745 58.480 46.975 61.140 ;
        RECT 46.710 55.680 47.010 58.480 ;
        RECT 46.745 53.140 46.975 55.680 ;
        RECT 49.035 54.530 49.265 61.140 ;
        RECT 50.375 61.030 50.605 61.140 ;
        RECT 50.340 59.630 50.640 61.030 ;
        RECT 49.000 53.130 49.300 54.530 ;
        RECT 50.375 53.140 50.605 59.630 ;
        RECT 52.665 58.480 52.895 61.140 ;
        RECT 52.630 55.680 52.930 58.480 ;
        RECT 52.665 53.140 52.895 55.680 ;
        RECT 54.955 54.530 55.185 61.140 ;
        RECT 57.245 58.480 57.475 61.140 ;
        RECT 59.535 61.030 59.765 61.140 ;
        RECT 59.500 59.630 59.800 61.030 ;
        RECT 57.210 55.680 57.510 58.480 ;
        RECT 54.920 53.130 55.220 54.530 ;
        RECT 57.245 53.140 57.475 55.680 ;
        RECT 59.535 53.140 59.765 59.630 ;
        RECT 61.825 58.480 62.055 61.140 ;
        RECT 61.790 55.680 62.090 58.480 ;
        RECT 61.825 53.140 62.055 55.680 ;
        RECT 64.115 54.530 64.345 61.140 ;
        RECT 66.405 58.480 66.635 61.140 ;
        RECT 68.695 61.030 68.925 61.140 ;
        RECT 70.035 61.030 70.265 61.140 ;
        RECT 68.660 59.630 68.960 61.030 ;
        RECT 70.000 59.630 70.300 61.030 ;
        RECT 66.370 55.680 66.670 58.480 ;
        RECT 64.080 53.130 64.380 54.530 ;
        RECT 66.405 53.140 66.635 55.680 ;
        RECT 68.695 53.140 68.925 59.630 ;
        RECT 70.035 53.140 70.265 59.630 ;
        RECT 72.325 58.480 72.555 61.140 ;
        RECT 72.290 55.680 72.590 58.480 ;
        RECT 72.325 53.140 72.555 55.680 ;
        RECT 74.615 54.530 74.845 61.140 ;
        RECT 76.905 58.480 77.135 61.140 ;
        RECT 79.195 61.030 79.425 61.140 ;
        RECT 79.160 59.630 79.460 61.030 ;
        RECT 76.870 55.680 77.170 58.480 ;
        RECT 74.580 53.130 74.880 54.530 ;
        RECT 76.905 53.140 77.135 55.680 ;
        RECT 79.195 53.140 79.425 59.630 ;
        RECT 81.485 58.480 81.715 61.140 ;
        RECT 81.450 55.680 81.750 58.480 ;
        RECT 81.485 53.140 81.715 55.680 ;
        RECT 83.775 54.530 84.005 61.140 ;
        RECT 86.065 58.480 86.295 61.140 ;
        RECT 88.355 61.030 88.585 61.140 ;
        RECT 88.320 59.630 88.620 61.030 ;
        RECT 86.030 55.680 86.330 58.480 ;
        RECT 83.740 53.130 84.040 54.530 ;
        RECT 86.065 53.140 86.295 55.680 ;
        RECT 88.355 53.140 88.585 59.630 ;
        RECT 89.695 54.530 89.925 61.140 ;
        RECT 91.985 58.480 92.215 61.140 ;
        RECT 94.275 61.030 94.505 61.140 ;
        RECT 94.240 59.630 94.540 61.030 ;
        RECT 91.950 55.680 92.250 58.480 ;
        RECT 89.660 53.130 89.960 54.530 ;
        RECT 91.985 53.140 92.215 55.680 ;
        RECT 94.275 53.140 94.505 59.630 ;
        RECT 96.565 58.480 96.795 61.140 ;
        RECT 96.530 55.680 96.830 58.480 ;
        RECT 96.565 53.140 96.795 55.680 ;
        RECT 98.855 54.530 99.085 61.140 ;
        RECT 101.145 58.480 101.375 61.140 ;
        RECT 103.435 61.030 103.665 61.140 ;
        RECT 103.400 59.630 103.700 61.030 ;
        RECT 101.110 55.680 101.410 58.480 ;
        RECT 98.820 53.130 99.120 54.530 ;
        RECT 101.145 53.140 101.375 55.680 ;
        RECT 103.435 53.140 103.665 59.630 ;
        RECT 105.725 58.480 105.955 61.140 ;
        RECT 105.690 55.680 105.990 58.480 ;
        RECT 105.725 53.140 105.955 55.680 ;
        RECT 108.015 54.530 108.245 61.140 ;
        RECT 107.980 53.130 108.280 54.530 ;
        RECT 109.355 52.935 109.585 61.345 ;
        RECT 111.645 52.935 111.875 61.345 ;
        RECT 113.935 52.935 114.165 61.345 ;
        RECT 116.225 52.935 116.455 61.345 ;
        RECT 118.515 52.935 118.745 61.345 ;
        RECT 120.805 52.935 121.035 61.345 ;
        RECT 123.095 52.935 123.325 61.345 ;
        RECT 125.385 52.935 125.615 61.345 ;
        RECT 127.675 52.935 127.905 61.345 ;
        RECT 11.055 51.325 29.605 52.935 ;
        RECT 30.995 52.705 32.955 52.935 ;
        RECT 33.285 52.345 35.245 52.935 ;
        RECT 35.575 52.345 37.535 52.935 ;
        RECT 37.865 52.705 39.825 52.935 ;
        RECT 40.155 52.705 42.115 52.935 ;
        RECT 42.445 52.345 44.405 52.935 ;
        RECT 44.735 52.345 46.695 52.935 ;
        RECT 47.025 52.705 48.985 52.935 ;
        RECT 50.655 52.345 52.615 52.935 ;
        RECT 52.945 52.705 54.905 52.935 ;
        RECT 55.235 52.705 57.195 52.935 ;
        RECT 57.525 52.345 59.485 52.935 ;
        RECT 59.815 52.345 61.775 52.935 ;
        RECT 62.105 52.705 64.065 52.935 ;
        RECT 64.395 52.705 66.355 52.935 ;
        RECT 66.685 52.345 68.645 52.935 ;
        RECT 70.315 52.345 72.275 52.935 ;
        RECT 72.605 52.705 74.565 52.935 ;
        RECT 74.895 52.705 76.855 52.935 ;
        RECT 77.185 52.345 79.145 52.935 ;
        RECT 79.475 52.345 81.435 52.935 ;
        RECT 81.765 52.705 83.725 52.935 ;
        RECT 84.055 52.705 86.015 52.935 ;
        RECT 86.345 52.345 88.305 52.935 ;
        RECT 89.975 52.705 91.935 52.935 ;
        RECT 92.265 52.345 94.225 52.935 ;
        RECT 94.555 52.345 96.515 52.935 ;
        RECT 96.845 52.705 98.805 52.935 ;
        RECT 99.135 52.705 101.095 52.935 ;
        RECT 101.425 52.345 103.385 52.935 ;
        RECT 103.715 52.345 105.675 52.935 ;
        RECT 106.005 52.705 107.965 52.935 ;
        RECT 30.995 51.325 32.955 51.555 ;
        RECT 33.285 51.325 35.245 51.555 ;
        RECT 35.575 51.325 37.535 51.555 ;
        RECT 37.865 51.325 39.825 51.555 ;
        RECT 40.155 51.325 42.115 51.555 ;
        RECT 42.445 51.325 44.405 51.555 ;
        RECT 44.735 51.325 46.695 51.555 ;
        RECT 47.025 51.325 48.985 51.555 ;
        RECT 50.655 51.325 52.615 51.555 ;
        RECT 52.945 51.325 54.905 51.555 ;
        RECT 55.235 51.325 57.195 51.555 ;
        RECT 57.525 51.325 59.485 51.555 ;
        RECT 59.815 51.325 61.775 51.555 ;
        RECT 62.105 51.325 64.065 51.555 ;
        RECT 64.395 51.325 66.355 51.555 ;
        RECT 66.685 51.325 68.645 51.555 ;
        RECT 70.315 51.325 72.275 51.555 ;
        RECT 72.605 51.325 74.565 51.555 ;
        RECT 74.895 51.325 76.855 51.555 ;
        RECT 77.185 51.325 79.145 51.555 ;
        RECT 79.475 51.325 81.435 51.555 ;
        RECT 81.765 51.325 83.725 51.555 ;
        RECT 84.055 51.325 86.015 51.555 ;
        RECT 86.345 51.325 88.305 51.555 ;
        RECT 89.975 51.325 91.935 51.555 ;
        RECT 92.265 51.325 94.225 51.555 ;
        RECT 94.555 51.325 96.515 51.555 ;
        RECT 96.845 51.325 98.805 51.555 ;
        RECT 99.135 51.325 101.095 51.555 ;
        RECT 101.425 51.325 103.385 51.555 ;
        RECT 103.715 51.325 105.675 51.555 ;
        RECT 106.005 51.325 107.965 51.555 ;
        RECT 109.355 51.325 127.905 52.935 ;
        RECT 11.055 42.915 11.285 51.325 ;
        RECT 13.345 42.915 13.575 51.325 ;
        RECT 15.635 42.915 15.865 51.325 ;
        RECT 17.925 42.915 18.155 51.325 ;
        RECT 20.215 42.915 20.445 51.325 ;
        RECT 22.505 42.915 22.735 51.325 ;
        RECT 24.795 42.915 25.025 51.325 ;
        RECT 27.085 42.915 27.315 51.325 ;
        RECT 29.375 42.915 29.605 51.325 ;
        RECT 11.055 42.225 29.605 42.915 ;
        RECT 30.715 42.915 30.945 51.120 ;
        RECT 33.005 42.915 33.235 51.120 ;
        RECT 35.295 42.915 35.525 51.120 ;
        RECT 37.585 42.915 37.815 51.120 ;
        RECT 39.875 42.915 40.105 51.120 ;
        RECT 42.165 42.915 42.395 51.120 ;
        RECT 44.455 42.915 44.685 51.120 ;
        RECT 46.745 42.915 46.975 51.120 ;
        RECT 49.035 42.915 49.265 51.120 ;
        RECT 30.715 42.225 49.265 42.915 ;
        RECT 50.375 42.915 50.605 51.120 ;
        RECT 52.665 42.915 52.895 51.120 ;
        RECT 54.955 42.915 55.185 51.120 ;
        RECT 57.245 42.915 57.475 51.120 ;
        RECT 59.535 42.915 59.765 51.120 ;
        RECT 61.825 42.915 62.055 51.120 ;
        RECT 64.115 42.915 64.345 51.120 ;
        RECT 66.405 42.915 66.635 51.120 ;
        RECT 68.695 42.915 68.925 51.120 ;
        RECT 50.375 42.225 68.925 42.915 ;
        RECT 70.035 42.915 70.265 51.120 ;
        RECT 72.325 42.915 72.555 51.120 ;
        RECT 74.615 42.915 74.845 51.120 ;
        RECT 76.905 42.915 77.135 51.120 ;
        RECT 79.195 42.915 79.425 51.120 ;
        RECT 81.485 42.915 81.715 51.120 ;
        RECT 83.775 42.915 84.005 51.120 ;
        RECT 86.065 42.915 86.295 51.120 ;
        RECT 88.355 42.915 88.585 51.120 ;
        RECT 70.035 42.225 88.585 42.915 ;
        RECT 89.695 42.915 89.925 51.120 ;
        RECT 91.985 42.915 92.215 51.120 ;
        RECT 94.275 42.915 94.505 51.120 ;
        RECT 96.565 42.915 96.795 51.120 ;
        RECT 98.855 42.915 99.085 51.120 ;
        RECT 101.145 42.915 101.375 51.120 ;
        RECT 103.435 42.915 103.665 51.120 ;
        RECT 105.725 42.915 105.955 51.120 ;
        RECT 108.015 42.915 108.245 51.120 ;
        RECT 89.695 42.225 108.245 42.915 ;
        RECT 109.355 42.915 109.585 51.325 ;
        RECT 111.645 42.915 111.875 51.325 ;
        RECT 113.935 42.915 114.165 51.325 ;
        RECT 116.225 42.915 116.455 51.325 ;
        RECT 118.515 42.915 118.745 51.325 ;
        RECT 120.805 42.915 121.035 51.325 ;
        RECT 123.095 42.915 123.325 51.325 ;
        RECT 125.385 42.915 125.615 51.325 ;
        RECT 127.675 42.915 127.905 51.325 ;
        RECT 109.355 42.225 127.905 42.915 ;
        RECT 128.345 42.225 135.710 102.115 ;
        RECT 136.295 100.155 138.400 101.915 ;
        RECT 136.295 97.815 138.400 99.575 ;
        RECT 136.295 95.475 138.400 97.235 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 141.695 93.725 142.995 108.925 ;
        RECT 149.570 107.765 155.900 137.690 ;
        RECT 234.845 109.385 235.165 109.445 ;
        RECT 263.365 109.385 263.685 109.445 ;
        RECT 234.845 109.245 263.685 109.385 ;
        RECT 234.845 109.185 235.165 109.245 ;
        RECT 263.365 109.185 263.685 109.245 ;
        RECT 232.085 109.045 232.405 109.105 ;
        RECT 253.245 109.045 253.565 109.105 ;
        RECT 232.085 108.905 253.565 109.045 ;
        RECT 232.085 108.845 232.405 108.905 ;
        RECT 253.245 108.845 253.565 108.905 ;
        RECT 238.985 108.705 239.305 108.765 ;
        RECT 259.685 108.705 260.005 108.765 ;
        RECT 238.985 108.565 260.005 108.705 ;
        RECT 238.985 108.505 239.305 108.565 ;
        RECT 259.685 108.505 260.005 108.565 ;
        RECT 209.085 108.365 209.405 108.425 ;
        RECT 254.625 108.365 254.945 108.425 ;
        RECT 209.085 108.225 254.945 108.365 ;
        RECT 209.085 108.165 209.405 108.225 ;
        RECT 254.625 108.165 254.945 108.225 ;
        RECT 221.965 108.025 222.285 108.085 ;
        RECT 240.825 108.025 241.145 108.085 ;
        RECT 221.965 107.885 241.145 108.025 ;
        RECT 221.965 107.825 222.285 107.885 ;
        RECT 240.825 107.825 241.145 107.885 ;
        RECT 248.645 108.025 248.965 108.085 ;
        RECT 261.525 108.025 261.845 108.085 ;
        RECT 248.645 107.885 261.845 108.025 ;
        RECT 248.645 107.825 248.965 107.885 ;
        RECT 261.525 107.825 261.845 107.885 ;
        RECT 146.290 104.835 155.900 107.765 ;
        RECT 171.825 107.685 172.145 107.745 ;
        RECT 184.705 107.685 185.025 107.745 ;
        RECT 171.825 107.545 185.025 107.685 ;
        RECT 171.825 107.485 172.145 107.545 ;
        RECT 184.705 107.485 185.025 107.545 ;
        RECT 252.785 107.685 253.105 107.745 ;
        RECT 261.985 107.685 262.305 107.745 ;
        RECT 252.785 107.545 262.305 107.685 ;
        RECT 252.785 107.485 253.105 107.545 ;
        RECT 261.985 107.485 262.305 107.545 ;
        RECT 272.105 107.685 272.425 107.745 ;
        RECT 282.685 107.685 283.005 107.745 ;
        RECT 272.105 107.545 283.005 107.685 ;
        RECT 272.105 107.485 272.425 107.545 ;
        RECT 282.685 107.485 283.005 107.545 ;
        RECT 172.285 107.345 172.605 107.405 ;
        RECT 229.325 107.345 229.645 107.405 ;
        RECT 257.845 107.345 258.165 107.405 ;
        RECT 172.285 107.205 184.935 107.345 ;
        RECT 172.285 107.145 172.605 107.205 ;
        RECT 184.795 107.065 184.935 107.205 ;
        RECT 229.325 107.205 258.165 107.345 ;
        RECT 229.325 107.145 229.645 107.205 ;
        RECT 257.845 107.145 258.165 107.205 ;
        RECT 258.305 107.345 258.625 107.405 ;
        RECT 276.705 107.345 277.025 107.405 ;
        RECT 258.305 107.205 277.025 107.345 ;
        RECT 258.305 107.145 258.625 107.205 ;
        RECT 276.705 107.145 277.025 107.205 ;
        RECT 168.145 107.005 168.465 107.065 ;
        RECT 177.805 107.005 178.125 107.065 ;
        RECT 168.145 106.865 178.125 107.005 ;
        RECT 168.145 106.805 168.465 106.865 ;
        RECT 177.805 106.805 178.125 106.865 ;
        RECT 184.705 106.805 185.025 107.065 ;
        RECT 204.025 107.005 204.345 107.065 ;
        RECT 210.005 107.005 210.325 107.065 ;
        RECT 204.025 106.865 210.325 107.005 ;
        RECT 204.025 106.805 204.345 106.865 ;
        RECT 210.005 106.805 210.325 106.865 ;
        RECT 244.505 107.005 244.825 107.065 ;
        RECT 264.285 107.005 264.605 107.065 ;
        RECT 244.505 106.865 264.605 107.005 ;
        RECT 244.505 106.805 244.825 106.865 ;
        RECT 264.285 106.805 264.605 106.865 ;
        RECT 279.005 107.005 279.325 107.065 ;
        RECT 304.765 107.005 305.085 107.065 ;
        RECT 279.005 106.865 305.085 107.005 ;
        RECT 279.005 106.805 279.325 106.865 ;
        RECT 304.765 106.805 305.085 106.865 ;
        RECT 162.095 106.185 311.135 106.665 ;
        RECT 164.480 105.985 164.770 106.030 ;
        RECT 173.205 105.985 173.525 106.045 ;
        RECT 164.480 105.845 173.525 105.985 ;
        RECT 164.480 105.800 164.770 105.845 ;
        RECT 173.205 105.785 173.525 105.845 ;
        RECT 174.140 105.985 174.430 106.030 ;
        RECT 174.140 105.845 180.335 105.985 ;
        RECT 174.140 105.800 174.430 105.845 ;
        RECT 173.665 105.645 173.985 105.705 ;
        RECT 173.665 105.505 177.115 105.645 ;
        RECT 173.665 105.445 173.985 105.505 ;
        RECT 176.975 105.365 177.115 105.505 ;
        RECT 164.465 105.305 164.785 105.365 ;
        RECT 165.400 105.305 165.690 105.350 ;
        RECT 164.465 105.165 165.690 105.305 ;
        RECT 164.465 105.105 164.785 105.165 ;
        RECT 165.400 105.120 165.690 105.165 ;
        RECT 166.765 105.305 167.085 105.365 ;
        RECT 167.240 105.305 167.530 105.350 ;
        RECT 166.765 105.165 167.530 105.305 ;
        RECT 166.765 105.105 167.085 105.165 ;
        RECT 167.240 105.120 167.530 105.165 ;
        RECT 169.065 105.105 169.385 105.365 ;
        RECT 170.920 105.305 171.210 105.350 ;
        RECT 172.285 105.305 172.605 105.365 ;
        RECT 170.920 105.165 172.605 105.305 ;
        RECT 170.920 105.120 171.210 105.165 ;
        RECT 172.285 105.105 172.605 105.165 ;
        RECT 172.745 105.105 173.065 105.365 ;
        RECT 173.220 105.305 173.510 105.350 ;
        RECT 174.585 105.305 174.905 105.365 ;
        RECT 173.220 105.165 174.905 105.305 ;
        RECT 173.220 105.120 173.510 105.165 ;
        RECT 174.585 105.105 174.905 105.165 ;
        RECT 175.045 105.305 175.365 105.365 ;
        RECT 176.885 105.305 177.205 105.365 ;
        RECT 177.360 105.305 177.650 105.350 ;
        RECT 175.045 105.165 176.655 105.305 ;
        RECT 175.045 105.105 175.365 105.165 ;
        RECT 175.505 104.965 175.825 105.025 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 146.290 101.325 148.395 103.085 ;
        RECT 146.290 98.985 148.395 100.745 ;
        RECT 146.290 96.645 148.395 98.405 ;
        RECT 146.290 94.305 148.395 96.065 ;
        RECT 136.295 91.965 138.400 93.725 ;
        RECT 141.695 93.135 148.395 93.725 ;
        RECT 146.290 91.965 148.395 92.555 ;
        RECT 136.295 90.795 143.395 91.385 ;
        RECT 136.295 89.625 138.400 90.215 ;
        RECT 146.290 89.625 148.395 91.385 ;
        RECT 136.295 87.285 138.400 89.045 ;
        RECT 146.290 88.455 148.395 89.045 ;
        RECT 146.290 87.285 148.395 87.875 ;
        RECT 136.295 86.115 138.400 86.705 ;
        RECT 136.295 84.945 138.400 85.535 ;
        RECT 146.290 84.945 148.395 86.705 ;
        RECT 136.295 82.605 138.400 84.365 ;
        RECT 146.290 83.775 148.395 84.365 ;
        RECT 146.290 82.605 148.395 83.195 ;
        RECT 136.295 81.435 141.260 82.025 ;
        RECT 143.790 81.435 148.395 82.025 ;
        RECT 136.295 80.265 138.400 80.855 ;
        RECT 136.295 79.095 138.400 79.685 ;
        RECT 136.295 76.755 138.400 78.515 ;
        RECT 136.295 75.585 138.400 76.175 ;
        RECT 136.295 74.415 138.400 75.005 ;
        RECT 136.295 72.075 138.400 73.835 ;
        RECT 136.295 70.905 138.400 71.495 ;
        RECT 136.295 69.735 138.400 70.325 ;
        RECT 136.295 67.395 138.400 69.155 ;
        RECT 136.295 66.225 138.400 66.815 ;
        RECT 136.295 65.055 138.400 65.645 ;
        RECT 136.295 62.715 138.400 64.475 ;
        RECT 143.790 62.135 145.190 81.435 ;
        RECT 146.290 79.095 148.395 80.855 ;
        RECT 146.290 77.925 148.395 78.515 ;
        RECT 146.290 76.755 148.395 77.345 ;
        RECT 146.290 74.415 148.395 76.175 ;
        RECT 146.290 73.245 148.395 73.835 ;
        RECT 146.290 72.075 148.395 72.665 ;
        RECT 146.290 69.735 148.395 71.495 ;
        RECT 146.290 68.565 148.395 69.155 ;
        RECT 146.290 67.395 148.395 67.985 ;
        RECT 146.290 65.055 148.395 66.815 ;
        RECT 146.290 63.885 148.395 64.475 ;
        RECT 146.290 62.715 148.395 63.305 ;
        RECT 136.295 61.545 140.910 62.135 ;
        RECT 143.790 61.545 148.395 62.135 ;
        RECT 136.295 60.375 138.400 60.965 ;
        RECT 136.295 59.205 138.400 59.795 ;
        RECT 136.295 56.865 138.400 58.625 ;
        RECT 136.295 55.695 138.400 56.285 ;
        RECT 136.295 54.525 138.400 55.115 ;
        RECT 136.295 52.185 138.400 53.945 ;
        RECT 136.295 51.015 138.400 51.605 ;
        RECT 136.295 49.845 138.400 50.435 ;
        RECT 136.295 47.505 138.400 49.265 ;
        RECT 136.295 46.335 138.400 46.925 ;
        RECT 136.295 45.165 138.400 45.755 ;
        RECT 136.295 42.825 138.400 44.585 ;
        RECT 139.510 42.245 140.910 61.545 ;
        RECT 146.290 59.205 148.395 60.965 ;
        RECT 146.290 58.035 148.395 58.625 ;
        RECT 146.290 56.865 148.395 57.455 ;
        RECT 146.290 54.525 148.395 56.285 ;
        RECT 146.290 53.355 148.395 53.945 ;
        RECT 146.290 52.185 148.395 52.775 ;
        RECT 146.290 49.845 148.395 51.605 ;
        RECT 146.290 48.675 148.395 49.265 ;
        RECT 146.290 47.505 148.395 48.095 ;
        RECT 146.290 45.165 148.395 46.925 ;
        RECT 146.290 43.995 148.395 44.585 ;
        RECT 146.290 42.825 148.395 43.415 ;
        RECT 4.100 41.635 135.710 42.225 ;
        RECT 136.295 41.655 140.910 42.245 ;
        RECT 143.435 41.655 148.395 42.245 ;
        RECT 4.100 4.900 4.900 41.635 ;
        RECT 7.065 39.040 130.565 39.630 ;
        RECT 7.065 36.430 10.615 39.040 ;
        RECT 8.665 9.480 10.615 36.430 ;
        RECT 11.115 38.350 20.505 38.580 ;
        RECT 22.015 38.350 30.845 38.650 ;
        RECT 32.635 38.350 41.465 38.650 ;
        RECT 43.255 38.350 52.085 38.650 ;
        RECT 53.875 38.350 62.705 38.650 ;
        RECT 64.215 38.350 73.605 38.580 ;
        RECT 11.115 34.890 11.345 38.350 ;
        RECT 13.405 34.890 13.635 38.190 ;
        RECT 15.695 34.890 15.925 38.350 ;
        RECT 17.985 34.890 18.215 38.190 ;
        RECT 20.275 34.890 20.505 38.350 ;
        RECT 11.020 33.490 11.345 34.890 ;
        RECT 13.370 33.490 13.670 34.890 ;
        RECT 15.660 33.490 15.960 34.890 ;
        RECT 17.950 33.490 18.250 34.890 ;
        RECT 20.240 33.490 20.540 34.890 ;
        RECT 11.115 30.030 11.345 33.490 ;
        RECT 13.405 30.190 13.635 33.490 ;
        RECT 15.695 30.030 15.925 33.490 ;
        RECT 17.985 30.190 18.215 33.490 ;
        RECT 20.275 30.030 20.505 33.490 ;
        RECT 21.735 32.890 21.965 38.190 ;
        RECT 24.025 34.890 24.255 38.190 ;
        RECT 26.315 36.890 26.545 38.190 ;
        RECT 26.280 35.490 26.580 36.890 ;
        RECT 23.990 33.490 24.290 34.890 ;
        RECT 21.700 31.490 22.000 32.890 ;
        RECT 21.735 30.190 21.965 31.490 ;
        RECT 24.025 30.190 24.255 33.490 ;
        RECT 26.315 30.190 26.545 35.490 ;
        RECT 28.605 34.890 28.835 38.190 ;
        RECT 28.570 33.490 28.870 34.890 ;
        RECT 28.605 30.190 28.835 33.490 ;
        RECT 30.895 32.890 31.125 38.190 ;
        RECT 32.355 36.890 32.585 38.190 ;
        RECT 32.320 35.490 32.620 36.890 ;
        RECT 30.860 31.490 31.160 32.890 ;
        RECT 30.895 30.190 31.125 31.490 ;
        RECT 32.355 30.190 32.585 35.490 ;
        RECT 34.645 34.890 34.875 38.190 ;
        RECT 34.610 33.490 34.910 34.890 ;
        RECT 34.645 30.190 34.875 33.490 ;
        RECT 36.935 32.890 37.165 38.190 ;
        RECT 39.225 34.890 39.455 38.190 ;
        RECT 41.515 36.890 41.745 38.190 ;
        RECT 41.480 35.490 41.780 36.890 ;
        RECT 39.190 33.490 39.490 34.890 ;
        RECT 36.900 31.490 37.200 32.890 ;
        RECT 36.935 30.190 37.165 31.490 ;
        RECT 39.225 30.190 39.455 33.490 ;
        RECT 41.515 30.190 41.745 35.490 ;
        RECT 42.975 32.890 43.205 38.190 ;
        RECT 45.265 34.890 45.495 38.190 ;
        RECT 47.555 36.890 47.785 38.190 ;
        RECT 47.520 35.490 47.820 36.890 ;
        RECT 45.230 33.490 45.530 34.890 ;
        RECT 42.940 31.490 43.240 32.890 ;
        RECT 42.975 30.190 43.205 31.490 ;
        RECT 45.265 30.190 45.495 33.490 ;
        RECT 47.555 30.190 47.785 35.490 ;
        RECT 49.845 34.890 50.075 38.190 ;
        RECT 49.810 33.490 50.110 34.890 ;
        RECT 49.845 30.190 50.075 33.490 ;
        RECT 52.135 32.890 52.365 38.190 ;
        RECT 53.595 36.890 53.825 38.190 ;
        RECT 53.560 35.490 53.860 36.890 ;
        RECT 52.100 31.490 52.400 32.890 ;
        RECT 52.135 30.190 52.365 31.490 ;
        RECT 53.595 30.190 53.825 35.490 ;
        RECT 55.885 34.890 56.115 38.190 ;
        RECT 55.850 33.490 56.150 34.890 ;
        RECT 55.885 30.190 56.115 33.490 ;
        RECT 58.175 32.890 58.405 38.190 ;
        RECT 60.465 34.890 60.695 38.190 ;
        RECT 62.755 36.890 62.985 38.190 ;
        RECT 62.720 35.490 63.020 36.890 ;
        RECT 60.430 33.490 60.730 34.890 ;
        RECT 58.140 31.490 58.440 32.890 ;
        RECT 58.175 30.190 58.405 31.490 ;
        RECT 60.465 30.190 60.695 33.490 ;
        RECT 62.755 30.190 62.985 35.490 ;
        RECT 64.215 34.890 64.445 38.350 ;
        RECT 66.505 34.890 66.735 38.190 ;
        RECT 68.795 34.890 69.025 38.350 ;
        RECT 71.085 34.890 71.315 38.190 ;
        RECT 73.375 34.890 73.605 38.350 ;
        RECT 64.180 33.490 64.480 34.890 ;
        RECT 66.470 33.490 66.770 34.890 ;
        RECT 68.760 33.490 69.060 34.890 ;
        RECT 71.050 33.490 71.350 34.890 ;
        RECT 73.340 33.490 73.640 34.890 ;
        RECT 64.215 30.030 64.445 33.490 ;
        RECT 66.505 30.190 66.735 33.490 ;
        RECT 68.795 30.030 69.025 33.490 ;
        RECT 71.085 30.190 71.315 33.490 ;
        RECT 73.375 30.030 73.605 33.490 ;
        RECT 11.115 29.800 20.505 30.030 ;
        RECT 22.015 29.730 30.845 30.030 ;
        RECT 32.635 29.730 41.465 30.030 ;
        RECT 43.255 29.730 52.085 30.030 ;
        RECT 53.875 29.730 62.705 30.030 ;
        RECT 64.215 29.800 73.605 30.030 ;
        RECT 11.115 28.420 20.505 28.650 ;
        RECT 22.015 28.420 30.845 28.720 ;
        RECT 32.635 28.650 41.465 28.720 ;
        RECT 43.255 28.650 52.085 28.720 ;
        RECT 32.355 28.420 41.745 28.650 ;
        RECT 11.115 24.960 11.345 28.420 ;
        RECT 13.405 24.960 13.635 28.260 ;
        RECT 15.695 24.960 15.925 28.420 ;
        RECT 17.985 24.960 18.215 28.260 ;
        RECT 20.275 24.960 20.505 28.420 ;
        RECT 21.735 26.960 21.965 28.260 ;
        RECT 21.700 25.560 22.000 26.960 ;
        RECT 11.020 23.560 11.345 24.960 ;
        RECT 13.370 23.560 13.670 24.960 ;
        RECT 15.660 23.560 15.960 24.960 ;
        RECT 17.950 23.560 18.250 24.960 ;
        RECT 20.240 23.560 20.540 24.960 ;
        RECT 11.115 20.100 11.345 23.560 ;
        RECT 13.405 20.260 13.635 23.560 ;
        RECT 15.695 20.100 15.925 23.560 ;
        RECT 17.985 20.260 18.215 23.560 ;
        RECT 20.275 20.100 20.505 23.560 ;
        RECT 21.735 20.260 21.965 25.560 ;
        RECT 24.025 24.960 24.255 28.260 ;
        RECT 23.990 23.560 24.290 24.960 ;
        RECT 24.025 20.260 24.255 23.560 ;
        RECT 26.315 22.960 26.545 28.260 ;
        RECT 28.605 24.960 28.835 28.260 ;
        RECT 30.895 26.960 31.125 28.260 ;
        RECT 30.860 25.560 31.160 26.960 ;
        RECT 28.570 23.560 28.870 24.960 ;
        RECT 26.280 21.560 26.580 22.960 ;
        RECT 26.315 20.260 26.545 21.560 ;
        RECT 28.605 20.260 28.835 23.560 ;
        RECT 30.895 20.260 31.125 25.560 ;
        RECT 32.355 20.100 32.585 28.420 ;
        RECT 34.645 24.960 34.875 28.260 ;
        RECT 34.610 23.560 34.910 24.960 ;
        RECT 34.645 20.260 34.875 23.560 ;
        RECT 36.935 20.100 37.165 28.420 ;
        RECT 39.225 24.960 39.455 28.260 ;
        RECT 39.190 23.560 39.490 24.960 ;
        RECT 39.225 20.260 39.455 23.560 ;
        RECT 41.515 20.100 41.745 28.420 ;
        RECT 11.115 19.870 20.505 20.100 ;
        RECT 22.015 19.800 30.845 20.100 ;
        RECT 32.355 19.870 41.745 20.100 ;
        RECT 42.975 28.420 52.365 28.650 ;
        RECT 53.875 28.420 62.705 28.720 ;
        RECT 64.215 28.420 73.605 28.650 ;
        RECT 42.975 20.100 43.205 28.420 ;
        RECT 45.265 24.960 45.495 28.260 ;
        RECT 45.230 23.560 45.530 24.960 ;
        RECT 45.265 20.260 45.495 23.560 ;
        RECT 47.555 20.100 47.785 28.420 ;
        RECT 49.845 24.960 50.075 28.260 ;
        RECT 49.810 23.560 50.110 24.960 ;
        RECT 49.845 20.260 50.075 23.560 ;
        RECT 52.135 20.100 52.365 28.420 ;
        RECT 53.595 22.960 53.825 28.260 ;
        RECT 55.885 24.960 56.115 28.260 ;
        RECT 58.175 26.960 58.405 28.260 ;
        RECT 58.140 25.560 58.440 26.960 ;
        RECT 55.850 23.560 56.150 24.960 ;
        RECT 53.560 21.560 53.860 22.960 ;
        RECT 53.595 20.260 53.825 21.560 ;
        RECT 55.885 20.260 56.115 23.560 ;
        RECT 58.175 20.260 58.405 25.560 ;
        RECT 60.465 24.960 60.695 28.260 ;
        RECT 60.430 23.560 60.730 24.960 ;
        RECT 60.465 20.260 60.695 23.560 ;
        RECT 62.755 22.960 62.985 28.260 ;
        RECT 64.215 24.960 64.445 28.420 ;
        RECT 66.505 24.960 66.735 28.260 ;
        RECT 68.795 24.960 69.025 28.420 ;
        RECT 71.085 24.960 71.315 28.260 ;
        RECT 73.375 24.960 73.605 28.420 ;
        RECT 64.180 23.560 64.480 24.960 ;
        RECT 66.470 23.560 66.770 24.960 ;
        RECT 68.760 23.560 69.060 24.960 ;
        RECT 71.050 23.560 71.350 24.960 ;
        RECT 73.340 23.560 73.640 24.960 ;
        RECT 62.720 21.560 63.020 22.960 ;
        RECT 62.755 20.260 62.985 21.560 ;
        RECT 64.215 20.100 64.445 23.560 ;
        RECT 66.505 20.260 66.735 23.560 ;
        RECT 68.795 20.100 69.025 23.560 ;
        RECT 71.085 20.260 71.315 23.560 ;
        RECT 73.375 20.100 73.605 23.560 ;
        RECT 42.975 19.870 52.365 20.100 ;
        RECT 32.635 19.800 41.465 19.870 ;
        RECT 43.255 19.800 52.085 19.870 ;
        RECT 53.875 19.800 62.705 20.100 ;
        RECT 64.215 19.870 73.605 20.100 ;
        RECT 11.115 18.490 20.505 18.720 ;
        RECT 22.015 18.490 30.845 18.790 ;
        RECT 32.635 18.490 41.465 18.790 ;
        RECT 43.255 18.490 52.085 18.790 ;
        RECT 53.875 18.490 62.705 18.790 ;
        RECT 64.215 18.490 73.605 18.720 ;
        RECT 11.115 15.030 11.345 18.490 ;
        RECT 13.405 15.030 13.635 18.330 ;
        RECT 15.695 15.030 15.925 18.490 ;
        RECT 17.985 15.030 18.215 18.330 ;
        RECT 20.275 15.030 20.505 18.490 ;
        RECT 11.020 13.630 11.345 15.030 ;
        RECT 13.370 13.630 13.670 15.030 ;
        RECT 15.660 13.630 15.960 15.030 ;
        RECT 17.950 13.630 18.250 15.030 ;
        RECT 20.240 13.630 20.540 15.030 ;
        RECT 11.115 10.170 11.345 13.630 ;
        RECT 13.405 10.330 13.635 13.630 ;
        RECT 15.695 10.170 15.925 13.630 ;
        RECT 17.985 10.330 18.215 13.630 ;
        RECT 20.275 10.170 20.505 13.630 ;
        RECT 21.735 13.030 21.965 18.330 ;
        RECT 24.025 15.030 24.255 18.330 ;
        RECT 26.315 17.030 26.545 18.330 ;
        RECT 26.280 15.630 26.580 17.030 ;
        RECT 23.990 13.630 24.290 15.030 ;
        RECT 21.700 11.630 22.000 13.030 ;
        RECT 21.735 10.330 21.965 11.630 ;
        RECT 24.025 10.330 24.255 13.630 ;
        RECT 26.315 10.330 26.545 15.630 ;
        RECT 28.605 15.030 28.835 18.330 ;
        RECT 28.570 13.630 28.870 15.030 ;
        RECT 28.605 10.330 28.835 13.630 ;
        RECT 30.895 13.030 31.125 18.330 ;
        RECT 32.355 17.030 32.585 18.330 ;
        RECT 32.320 15.630 32.620 17.030 ;
        RECT 30.860 11.630 31.160 13.030 ;
        RECT 30.895 10.330 31.125 11.630 ;
        RECT 32.355 10.330 32.585 15.630 ;
        RECT 34.645 15.030 34.875 18.330 ;
        RECT 34.610 13.630 34.910 15.030 ;
        RECT 34.645 10.330 34.875 13.630 ;
        RECT 36.935 13.030 37.165 18.330 ;
        RECT 39.225 15.030 39.455 18.330 ;
        RECT 41.515 17.030 41.745 18.330 ;
        RECT 41.480 15.630 41.780 17.030 ;
        RECT 39.190 13.630 39.490 15.030 ;
        RECT 36.900 11.630 37.200 13.030 ;
        RECT 36.935 10.330 37.165 11.630 ;
        RECT 39.225 10.330 39.455 13.630 ;
        RECT 41.515 10.330 41.745 15.630 ;
        RECT 42.975 13.030 43.205 18.330 ;
        RECT 45.265 15.030 45.495 18.330 ;
        RECT 47.555 17.030 47.785 18.330 ;
        RECT 47.520 15.630 47.820 17.030 ;
        RECT 45.230 13.630 45.530 15.030 ;
        RECT 42.940 11.630 43.240 13.030 ;
        RECT 42.975 10.330 43.205 11.630 ;
        RECT 45.265 10.330 45.495 13.630 ;
        RECT 47.555 10.330 47.785 15.630 ;
        RECT 49.845 15.030 50.075 18.330 ;
        RECT 49.810 13.630 50.110 15.030 ;
        RECT 49.845 10.330 50.075 13.630 ;
        RECT 52.135 13.030 52.365 18.330 ;
        RECT 53.595 17.030 53.825 18.330 ;
        RECT 53.560 15.630 53.860 17.030 ;
        RECT 52.100 11.630 52.400 13.030 ;
        RECT 52.135 10.330 52.365 11.630 ;
        RECT 53.595 10.330 53.825 15.630 ;
        RECT 55.885 15.030 56.115 18.330 ;
        RECT 55.850 13.630 56.150 15.030 ;
        RECT 55.885 10.330 56.115 13.630 ;
        RECT 58.175 13.030 58.405 18.330 ;
        RECT 60.465 15.030 60.695 18.330 ;
        RECT 62.755 17.030 62.985 18.330 ;
        RECT 62.720 15.630 63.020 17.030 ;
        RECT 60.430 13.630 60.730 15.030 ;
        RECT 58.140 11.630 58.440 13.030 ;
        RECT 58.175 10.330 58.405 11.630 ;
        RECT 60.465 10.330 60.695 13.630 ;
        RECT 62.755 10.330 62.985 15.630 ;
        RECT 64.215 15.030 64.445 18.490 ;
        RECT 66.505 15.030 66.735 18.330 ;
        RECT 68.795 15.030 69.025 18.490 ;
        RECT 71.085 15.030 71.315 18.330 ;
        RECT 73.375 15.030 73.605 18.490 ;
        RECT 64.180 13.630 64.480 15.030 ;
        RECT 66.470 13.630 66.770 15.030 ;
        RECT 68.760 13.630 69.060 15.030 ;
        RECT 71.050 13.630 71.350 15.030 ;
        RECT 73.340 13.630 73.640 15.030 ;
        RECT 64.215 10.170 64.445 13.630 ;
        RECT 66.505 10.330 66.735 13.630 ;
        RECT 68.795 10.170 69.025 13.630 ;
        RECT 71.085 10.330 71.315 13.630 ;
        RECT 73.375 10.170 73.605 13.630 ;
        RECT 11.115 9.940 20.505 10.170 ;
        RECT 22.015 9.870 30.845 10.170 ;
        RECT 32.635 9.870 41.465 10.170 ;
        RECT 43.255 9.870 52.085 10.170 ;
        RECT 53.875 9.870 62.705 10.170 ;
        RECT 64.215 9.940 73.605 10.170 ;
        RECT 74.105 9.480 80.255 39.040 ;
        RECT 81.035 38.350 82.995 38.580 ;
        RECT 83.325 38.350 85.285 38.580 ;
        RECT 87.075 38.350 89.035 38.700 ;
        RECT 89.365 38.350 91.325 38.700 ;
        RECT 93.115 38.350 97.365 38.700 ;
        RECT 99.155 38.350 101.115 38.700 ;
        RECT 101.445 38.350 103.405 38.700 ;
        RECT 105.195 38.350 107.155 38.700 ;
        RECT 107.485 38.350 109.445 38.700 ;
        RECT 111.235 38.350 115.485 38.700 ;
        RECT 117.275 38.350 119.235 38.700 ;
        RECT 119.565 38.350 121.525 38.700 ;
        RECT 123.315 38.350 125.275 38.580 ;
        RECT 125.605 38.350 127.565 38.580 ;
        RECT 80.755 30.190 80.985 38.190 ;
        RECT 83.045 30.190 83.275 38.190 ;
        RECT 85.335 30.190 85.565 38.190 ;
        RECT 86.795 35.995 87.025 38.190 ;
        RECT 86.560 35.295 87.260 35.995 ;
        RECT 86.795 30.190 87.025 35.295 ;
        RECT 89.085 34.495 89.315 38.190 ;
        RECT 91.375 35.995 91.605 38.190 ;
        RECT 92.835 37.495 93.065 38.190 ;
        RECT 92.600 36.795 93.300 37.495 ;
        RECT 91.140 35.295 91.840 35.995 ;
        RECT 88.850 33.795 89.550 34.495 ;
        RECT 89.085 30.190 89.315 33.795 ;
        RECT 91.375 30.190 91.605 35.295 ;
        RECT 92.835 30.190 93.065 36.795 ;
        RECT 95.125 30.190 95.355 38.350 ;
        RECT 97.415 37.495 97.645 38.190 ;
        RECT 97.180 36.795 97.880 37.495 ;
        RECT 97.415 30.190 97.645 36.795 ;
        RECT 98.875 31.495 99.105 38.190 ;
        RECT 101.165 32.995 101.395 38.190 ;
        RECT 100.930 32.295 101.630 32.995 ;
        RECT 98.640 30.795 99.340 31.495 ;
        RECT 98.875 30.190 99.105 30.795 ;
        RECT 101.165 30.190 101.395 32.295 ;
        RECT 103.455 31.495 103.685 38.190 ;
        RECT 104.915 31.495 105.145 38.190 ;
        RECT 107.205 32.995 107.435 38.190 ;
        RECT 106.970 32.295 107.670 32.995 ;
        RECT 103.220 30.795 103.920 31.495 ;
        RECT 104.680 30.795 105.380 31.495 ;
        RECT 103.455 30.190 103.685 30.795 ;
        RECT 104.915 30.190 105.145 30.795 ;
        RECT 107.205 30.190 107.435 32.295 ;
        RECT 109.495 31.495 109.725 38.190 ;
        RECT 110.955 37.495 111.185 38.190 ;
        RECT 110.720 36.795 111.420 37.495 ;
        RECT 109.260 30.795 109.960 31.495 ;
        RECT 109.495 30.190 109.725 30.795 ;
        RECT 110.955 30.190 111.185 36.795 ;
        RECT 113.245 30.190 113.475 38.350 ;
        RECT 115.535 37.495 115.765 38.190 ;
        RECT 115.300 36.795 116.000 37.495 ;
        RECT 115.535 30.190 115.765 36.795 ;
        RECT 116.995 35.995 117.225 38.190 ;
        RECT 116.760 35.295 117.460 35.995 ;
        RECT 116.995 30.190 117.225 35.295 ;
        RECT 119.285 34.495 119.515 38.190 ;
        RECT 121.575 35.995 121.805 38.190 ;
        RECT 121.340 35.295 122.040 35.995 ;
        RECT 119.050 33.795 119.750 34.495 ;
        RECT 119.285 30.190 119.515 33.795 ;
        RECT 121.575 30.190 121.805 35.295 ;
        RECT 123.035 30.190 123.265 38.190 ;
        RECT 125.325 30.190 125.555 38.190 ;
        RECT 127.615 30.190 127.845 38.190 ;
        RECT 81.035 29.800 82.995 30.030 ;
        RECT 83.325 29.800 85.285 30.030 ;
        RECT 87.075 29.680 89.035 30.030 ;
        RECT 89.365 29.680 91.325 30.030 ;
        RECT 93.115 29.680 95.075 30.030 ;
        RECT 95.405 29.680 97.365 30.030 ;
        RECT 99.155 29.680 101.115 30.030 ;
        RECT 101.445 29.680 103.405 30.030 ;
        RECT 105.195 29.680 107.155 30.030 ;
        RECT 107.485 29.680 109.445 30.030 ;
        RECT 111.235 29.680 113.195 30.030 ;
        RECT 113.525 29.680 115.485 30.030 ;
        RECT 117.275 29.680 119.235 30.030 ;
        RECT 119.565 29.680 121.525 30.030 ;
        RECT 123.315 29.800 125.275 30.030 ;
        RECT 125.605 29.800 127.565 30.030 ;
        RECT 81.035 28.420 82.995 28.650 ;
        RECT 83.325 28.420 85.285 28.650 ;
        RECT 87.075 28.420 89.035 28.770 ;
        RECT 89.365 28.420 91.325 28.770 ;
        RECT 93.115 28.420 95.075 28.770 ;
        RECT 95.405 28.420 97.365 28.770 ;
        RECT 99.155 28.420 101.115 28.770 ;
        RECT 101.445 28.420 103.405 28.770 ;
        RECT 105.195 28.420 107.155 28.770 ;
        RECT 107.485 28.420 109.445 28.770 ;
        RECT 111.235 28.420 113.195 28.770 ;
        RECT 113.525 28.420 115.485 28.770 ;
        RECT 117.275 28.420 119.235 28.770 ;
        RECT 119.565 28.420 121.525 28.770 ;
        RECT 123.315 28.420 125.275 28.650 ;
        RECT 125.605 28.420 127.565 28.650 ;
        RECT 80.755 20.260 80.985 28.260 ;
        RECT 83.045 20.260 83.275 28.260 ;
        RECT 85.335 20.260 85.565 28.260 ;
        RECT 86.795 23.065 87.025 28.260 ;
        RECT 89.085 24.565 89.315 28.260 ;
        RECT 88.850 23.865 89.550 24.565 ;
        RECT 86.560 22.365 87.260 23.065 ;
        RECT 86.795 20.260 87.025 22.365 ;
        RECT 89.085 20.260 89.315 23.865 ;
        RECT 91.375 23.065 91.605 28.260 ;
        RECT 91.140 22.365 91.840 23.065 ;
        RECT 91.375 20.260 91.605 22.365 ;
        RECT 92.835 21.565 93.065 28.260 ;
        RECT 92.600 20.865 93.300 21.565 ;
        RECT 92.835 20.260 93.065 20.865 ;
        RECT 95.125 20.100 95.355 28.260 ;
        RECT 97.415 21.565 97.645 28.260 ;
        RECT 98.875 27.565 99.105 28.260 ;
        RECT 98.640 26.865 99.340 27.565 ;
        RECT 97.180 20.865 97.880 21.565 ;
        RECT 97.415 20.260 97.645 20.865 ;
        RECT 98.875 20.260 99.105 26.865 ;
        RECT 101.165 26.065 101.395 28.260 ;
        RECT 103.455 27.565 103.685 28.260 ;
        RECT 104.915 27.565 105.145 28.260 ;
        RECT 103.220 26.865 103.920 27.565 ;
        RECT 104.680 26.865 105.380 27.565 ;
        RECT 100.930 25.365 101.630 26.065 ;
        RECT 101.165 20.260 101.395 25.365 ;
        RECT 103.455 20.260 103.685 26.865 ;
        RECT 104.915 20.260 105.145 26.865 ;
        RECT 107.205 26.065 107.435 28.260 ;
        RECT 109.495 27.565 109.725 28.260 ;
        RECT 109.260 26.865 109.960 27.565 ;
        RECT 106.970 25.365 107.670 26.065 ;
        RECT 107.205 20.260 107.435 25.365 ;
        RECT 109.495 20.260 109.725 26.865 ;
        RECT 110.955 21.565 111.185 28.260 ;
        RECT 110.720 20.865 111.420 21.565 ;
        RECT 110.955 20.260 111.185 20.865 ;
        RECT 113.245 20.100 113.475 28.260 ;
        RECT 115.535 21.565 115.765 28.260 ;
        RECT 116.995 23.065 117.225 28.260 ;
        RECT 119.285 24.565 119.515 28.260 ;
        RECT 119.050 23.865 119.750 24.565 ;
        RECT 116.760 22.365 117.460 23.065 ;
        RECT 115.300 20.865 116.000 21.565 ;
        RECT 115.535 20.260 115.765 20.865 ;
        RECT 116.995 20.260 117.225 22.365 ;
        RECT 119.285 20.260 119.515 23.865 ;
        RECT 121.575 23.065 121.805 28.260 ;
        RECT 121.340 22.365 122.040 23.065 ;
        RECT 121.575 20.260 121.805 22.365 ;
        RECT 123.035 20.260 123.265 28.260 ;
        RECT 125.325 20.260 125.555 28.260 ;
        RECT 127.615 20.260 127.845 28.260 ;
        RECT 81.035 19.870 82.995 20.100 ;
        RECT 83.325 19.870 85.285 20.100 ;
        RECT 87.075 19.750 89.035 20.100 ;
        RECT 89.365 19.750 91.325 20.100 ;
        RECT 93.115 19.750 97.365 20.100 ;
        RECT 99.155 19.750 101.115 20.100 ;
        RECT 101.445 19.750 103.405 20.100 ;
        RECT 105.195 19.750 107.155 20.100 ;
        RECT 107.485 19.750 109.445 20.100 ;
        RECT 111.235 19.750 115.485 20.100 ;
        RECT 117.275 19.750 119.235 20.100 ;
        RECT 119.565 19.750 121.525 20.100 ;
        RECT 123.315 19.870 125.275 20.100 ;
        RECT 125.605 19.870 127.565 20.100 ;
        RECT 81.035 18.490 82.995 18.720 ;
        RECT 83.325 18.490 85.285 18.720 ;
        RECT 87.075 18.490 89.035 18.720 ;
        RECT 89.365 18.490 91.325 18.720 ;
        RECT 93.115 18.490 95.075 18.720 ;
        RECT 95.405 18.490 97.365 18.720 ;
        RECT 99.155 18.490 101.115 18.720 ;
        RECT 101.445 18.490 103.405 18.720 ;
        RECT 105.195 18.490 107.155 18.720 ;
        RECT 107.485 18.490 109.445 18.720 ;
        RECT 111.235 18.490 113.195 18.720 ;
        RECT 113.525 18.490 115.485 18.720 ;
        RECT 117.275 18.490 119.235 18.720 ;
        RECT 119.565 18.490 121.525 18.720 ;
        RECT 123.315 18.490 125.275 18.720 ;
        RECT 125.605 18.490 127.565 18.720 ;
        RECT 80.755 10.330 80.985 18.330 ;
        RECT 83.045 10.330 83.275 18.330 ;
        RECT 85.335 10.330 85.565 18.330 ;
        RECT 86.795 10.330 87.025 18.330 ;
        RECT 89.085 10.330 89.315 18.330 ;
        RECT 91.375 10.330 91.605 18.330 ;
        RECT 92.835 10.330 93.065 18.330 ;
        RECT 95.125 10.330 95.355 18.330 ;
        RECT 97.415 10.330 97.645 18.330 ;
        RECT 98.875 10.330 99.105 18.330 ;
        RECT 101.165 10.330 101.395 18.330 ;
        RECT 103.455 10.330 103.685 18.330 ;
        RECT 104.915 10.330 105.145 18.330 ;
        RECT 107.205 10.330 107.435 18.330 ;
        RECT 109.495 10.330 109.725 18.330 ;
        RECT 110.955 10.330 111.185 18.330 ;
        RECT 113.245 10.330 113.475 18.330 ;
        RECT 115.535 10.330 115.765 18.330 ;
        RECT 116.995 10.330 117.225 18.330 ;
        RECT 119.285 10.330 119.515 18.330 ;
        RECT 121.575 10.330 121.805 18.330 ;
        RECT 123.035 10.330 123.265 18.330 ;
        RECT 125.325 10.330 125.555 18.330 ;
        RECT 127.615 10.330 127.845 18.330 ;
        RECT 81.035 9.940 82.995 10.170 ;
        RECT 83.325 9.940 85.285 10.170 ;
        RECT 87.075 9.940 89.035 10.170 ;
        RECT 89.365 9.940 91.325 10.170 ;
        RECT 93.115 9.940 95.075 10.170 ;
        RECT 95.405 9.940 97.365 10.170 ;
        RECT 99.155 9.940 101.115 10.170 ;
        RECT 101.445 9.940 103.405 10.170 ;
        RECT 105.195 9.940 107.155 10.170 ;
        RECT 107.485 9.940 109.445 10.170 ;
        RECT 111.235 9.940 113.195 10.170 ;
        RECT 113.525 9.940 115.485 10.170 ;
        RECT 117.275 9.940 119.235 10.170 ;
        RECT 119.565 9.940 121.525 10.170 ;
        RECT 123.315 9.940 125.275 10.170 ;
        RECT 125.605 9.940 127.565 10.170 ;
        RECT 128.345 9.480 130.565 39.040 ;
        RECT 8.665 8.890 130.565 9.480 ;
        RECT 7.065 5.690 130.565 8.890 ;
        RECT 135.120 18.845 135.710 41.635 ;
        RECT 136.295 40.485 138.400 41.075 ;
        RECT 136.295 39.315 138.400 39.905 ;
        RECT 146.290 39.315 148.395 41.075 ;
        RECT 136.295 36.975 138.400 38.735 ;
        RECT 146.290 38.145 148.395 38.735 ;
        RECT 146.290 36.975 148.395 37.565 ;
        RECT 136.295 35.805 138.400 36.395 ;
        RECT 136.295 34.635 138.400 35.225 ;
        RECT 146.290 34.635 148.395 36.395 ;
        RECT 136.295 32.295 138.400 34.055 ;
        RECT 146.290 33.465 148.395 34.055 ;
        RECT 143.640 32.295 148.395 32.885 ;
        RECT 136.295 31.125 138.400 31.715 ;
        RECT 136.295 29.955 141.055 30.545 ;
        RECT 146.290 29.955 148.395 31.715 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 136.295 26.445 138.400 28.205 ;
        RECT 146.290 27.615 148.395 29.375 ;
        RECT 136.295 24.105 138.400 25.865 ;
        RECT 146.290 25.275 148.395 27.035 ;
        RECT 136.295 21.765 138.400 23.525 ;
        RECT 146.290 22.935 148.395 24.695 ;
        RECT 136.295 19.425 138.400 21.185 ;
        RECT 146.290 20.595 148.395 22.355 ;
        RECT 141.295 19.425 148.395 20.015 ;
        RECT 148.980 18.845 155.900 104.835 ;
        RECT 169.615 104.825 175.825 104.965 ;
        RECT 176.515 104.965 176.655 105.165 ;
        RECT 176.885 105.165 177.650 105.305 ;
        RECT 176.885 105.105 177.205 105.165 ;
        RECT 177.360 105.120 177.650 105.165 ;
        RECT 177.820 104.965 178.110 105.010 ;
        RECT 176.515 104.825 178.110 104.965 ;
        RECT 168.145 104.425 168.465 104.685 ;
        RECT 166.320 104.285 166.610 104.330 ;
        RECT 169.615 104.285 169.755 104.825 ;
        RECT 175.505 104.765 175.825 104.825 ;
        RECT 177.820 104.780 178.110 104.825 ;
        RECT 178.740 104.965 179.030 105.010 ;
        RECT 179.645 104.965 179.965 105.025 ;
        RECT 178.740 104.825 179.965 104.965 ;
        RECT 180.195 104.965 180.335 105.845 ;
        RECT 181.500 105.800 181.790 106.030 ;
        RECT 183.340 105.985 183.630 106.030 ;
        RECT 193.905 105.985 194.225 106.045 ;
        RECT 183.340 105.845 194.225 105.985 ;
        RECT 183.340 105.800 183.630 105.845 ;
        RECT 181.575 105.645 181.715 105.800 ;
        RECT 193.905 105.785 194.225 105.845 ;
        RECT 199.900 105.985 200.190 106.030 ;
        RECT 205.405 105.985 205.725 106.045 ;
        RECT 208.165 105.985 208.485 106.045 ;
        RECT 199.900 105.845 205.725 105.985 ;
        RECT 199.900 105.800 200.190 105.845 ;
        RECT 205.405 105.785 205.725 105.845 ;
        RECT 206.415 105.845 208.485 105.985 ;
        RECT 191.145 105.645 191.465 105.705 ;
        RECT 192.525 105.690 192.845 105.705 ;
        RECT 181.575 105.505 191.465 105.645 ;
        RECT 191.145 105.445 191.465 105.505 ;
        RECT 192.060 105.645 192.845 105.690 ;
        RECT 195.660 105.645 195.950 105.690 ;
        RECT 206.415 105.645 206.555 105.845 ;
        RECT 208.165 105.785 208.485 105.845 ;
        RECT 209.085 105.785 209.405 106.045 ;
        RECT 212.320 105.985 212.610 106.030 ;
        RECT 216.905 105.985 217.225 106.045 ;
        RECT 212.320 105.845 217.225 105.985 ;
        RECT 212.320 105.800 212.610 105.845 ;
        RECT 216.905 105.785 217.225 105.845 ;
        RECT 218.760 105.985 219.050 106.030 ;
        RECT 223.805 105.985 224.125 106.045 ;
        RECT 218.760 105.845 224.125 105.985 ;
        RECT 218.760 105.800 219.050 105.845 ;
        RECT 223.805 105.785 224.125 105.845 ;
        RECT 225.200 105.985 225.490 106.030 ;
        RECT 228.405 105.985 228.725 106.045 ;
        RECT 225.200 105.845 228.725 105.985 ;
        RECT 225.200 105.800 225.490 105.845 ;
        RECT 228.405 105.785 228.725 105.845 ;
        RECT 230.705 105.985 231.025 106.045 ;
        RECT 231.640 105.985 231.930 106.030 ;
        RECT 230.705 105.845 231.930 105.985 ;
        RECT 230.705 105.785 231.025 105.845 ;
        RECT 231.640 105.800 231.930 105.845 ;
        RECT 233.005 105.985 233.325 106.045 ;
        RECT 233.940 105.985 234.230 106.030 ;
        RECT 233.005 105.845 234.230 105.985 ;
        RECT 233.005 105.785 233.325 105.845 ;
        RECT 233.940 105.800 234.230 105.845 ;
        RECT 235.305 105.985 235.625 106.045 ;
        RECT 236.700 105.985 236.990 106.030 ;
        RECT 235.305 105.845 236.990 105.985 ;
        RECT 235.305 105.785 235.625 105.845 ;
        RECT 236.700 105.800 236.990 105.845 ;
        RECT 237.605 105.985 237.925 106.045 ;
        RECT 238.080 105.985 238.370 106.030 ;
        RECT 237.605 105.845 238.370 105.985 ;
        RECT 237.605 105.785 237.925 105.845 ;
        RECT 238.080 105.800 238.370 105.845 ;
        RECT 242.205 105.785 242.525 106.045 ;
        RECT 249.105 105.985 249.425 106.045 ;
        RECT 266.140 105.985 266.430 106.030 ;
        RECT 249.105 105.845 266.430 105.985 ;
        RECT 249.105 105.785 249.425 105.845 ;
        RECT 266.140 105.800 266.430 105.845 ;
        RECT 269.820 105.800 270.110 106.030 ;
        RECT 221.520 105.645 221.810 105.690 ;
        RECT 227.040 105.645 227.330 105.690 ;
        RECT 192.060 105.505 195.950 105.645 ;
        RECT 192.060 105.460 192.845 105.505 ;
        RECT 192.525 105.445 192.845 105.460 ;
        RECT 195.360 105.460 195.950 105.505 ;
        RECT 201.355 105.505 206.555 105.645 ;
        RECT 215.155 105.505 218.515 105.645 ;
        RECT 180.565 105.105 180.885 105.365 ;
        RECT 182.420 105.305 182.710 105.350 ;
        RECT 183.325 105.305 183.645 105.365 ;
        RECT 182.420 105.165 183.645 105.305 ;
        RECT 182.420 105.120 182.710 105.165 ;
        RECT 183.325 105.105 183.645 105.165 ;
        RECT 188.865 105.305 189.155 105.350 ;
        RECT 190.700 105.305 190.990 105.350 ;
        RECT 194.280 105.305 194.570 105.350 ;
        RECT 188.865 105.165 194.570 105.305 ;
        RECT 188.865 105.120 189.155 105.165 ;
        RECT 190.700 105.120 190.990 105.165 ;
        RECT 194.280 105.120 194.570 105.165 ;
        RECT 195.360 105.145 195.650 105.460 ;
        RECT 198.965 105.105 199.285 105.365 ;
        RECT 201.355 105.350 201.495 105.505 ;
        RECT 201.280 105.120 201.570 105.350 ;
        RECT 202.185 105.305 202.505 105.365 ;
        RECT 203.120 105.305 203.410 105.350 ;
        RECT 205.865 105.305 206.185 105.365 ;
        RECT 206.340 105.305 206.630 105.350 ;
        RECT 202.185 105.165 203.410 105.305 ;
        RECT 186.545 104.965 186.865 105.025 ;
        RECT 180.195 104.825 186.865 104.965 ;
        RECT 178.740 104.780 179.030 104.825 ;
        RECT 179.645 104.765 179.965 104.825 ;
        RECT 186.545 104.765 186.865 104.825 ;
        RECT 187.480 104.780 187.770 105.010 ;
        RECT 170.000 104.625 170.290 104.670 ;
        RECT 180.105 104.625 180.425 104.685 ;
        RECT 170.000 104.485 180.425 104.625 ;
        RECT 170.000 104.440 170.290 104.485 ;
        RECT 180.105 104.425 180.425 104.485 ;
        RECT 166.320 104.145 169.755 104.285 ;
        RECT 166.320 104.100 166.610 104.145 ;
        RECT 171.825 104.085 172.145 104.345 ;
        RECT 175.505 104.085 175.825 104.345 ;
        RECT 184.245 104.085 184.565 104.345 ;
        RECT 187.555 104.285 187.695 104.780 ;
        RECT 188.385 104.765 188.705 105.025 ;
        RECT 189.765 104.765 190.085 105.025 ;
        RECT 201.355 104.965 201.495 105.120 ;
        RECT 202.185 105.105 202.505 105.165 ;
        RECT 203.120 105.120 203.410 105.165 ;
        RECT 204.575 105.165 205.635 105.305 ;
        RECT 204.575 104.965 204.715 105.165 ;
        RECT 197.215 104.825 201.495 104.965 ;
        RECT 202.275 104.825 204.715 104.965 ;
        RECT 189.270 104.625 189.560 104.670 ;
        RECT 191.160 104.625 191.450 104.670 ;
        RECT 194.280 104.625 194.570 104.670 ;
        RECT 189.270 104.485 194.570 104.625 ;
        RECT 189.270 104.440 189.560 104.485 ;
        RECT 191.160 104.440 191.450 104.485 ;
        RECT 194.280 104.440 194.570 104.485 ;
        RECT 197.215 104.330 197.355 104.825 ;
        RECT 202.275 104.670 202.415 104.825 ;
        RECT 202.200 104.440 202.490 104.670 ;
        RECT 204.025 104.425 204.345 104.685 ;
        RECT 205.495 104.625 205.635 105.165 ;
        RECT 205.865 105.165 206.630 105.305 ;
        RECT 205.865 105.105 206.185 105.165 ;
        RECT 206.340 105.120 206.630 105.165 ;
        RECT 208.625 105.105 208.945 105.365 ;
        RECT 213.225 105.105 213.545 105.365 ;
        RECT 210.020 104.965 210.310 105.010 ;
        RECT 215.155 104.965 215.295 105.505 ;
        RECT 218.375 105.365 218.515 105.505 ;
        RECT 221.520 105.505 227.330 105.645 ;
        RECT 221.520 105.460 221.810 105.505 ;
        RECT 227.040 105.460 227.330 105.505 ;
        RECT 230.245 105.645 230.565 105.705 ;
        RECT 242.295 105.645 242.435 105.785 ;
        RECT 253.705 105.645 254.025 105.705 ;
        RECT 269.895 105.645 270.035 105.800 ;
        RECT 276.705 105.785 277.025 106.045 ;
        RECT 291.900 105.985 292.190 106.030 ;
        RECT 279.555 105.845 292.190 105.985 ;
        RECT 230.245 105.505 235.995 105.645 ;
        RECT 242.295 105.505 252.555 105.645 ;
        RECT 230.245 105.445 230.565 105.505 ;
        RECT 215.540 105.305 215.830 105.350 ;
        RECT 216.905 105.305 217.225 105.365 ;
        RECT 215.540 105.165 217.225 105.305 ;
        RECT 215.540 105.120 215.830 105.165 ;
        RECT 216.905 105.105 217.225 105.165 ;
        RECT 217.365 105.105 217.685 105.365 ;
        RECT 217.825 105.105 218.145 105.365 ;
        RECT 218.285 105.305 218.605 105.365 ;
        RECT 226.120 105.305 226.410 105.350 ;
        RECT 232.085 105.305 232.405 105.365 ;
        RECT 218.285 105.165 222.655 105.305 ;
        RECT 218.285 105.105 218.605 105.165 ;
        RECT 221.505 104.965 221.825 105.025 ;
        RECT 210.020 104.825 215.295 104.965 ;
        RECT 216.995 104.825 221.825 104.965 ;
        RECT 210.020 104.780 210.310 104.825 ;
        RECT 207.705 104.625 208.025 104.685 ;
        RECT 205.495 104.485 208.025 104.625 ;
        RECT 207.705 104.425 208.025 104.485 ;
        RECT 216.460 104.625 216.750 104.670 ;
        RECT 216.995 104.625 217.135 104.825 ;
        RECT 221.505 104.765 221.825 104.825 ;
        RECT 221.965 104.765 222.285 105.025 ;
        RECT 222.515 105.010 222.655 105.165 ;
        RECT 226.120 105.165 232.405 105.305 ;
        RECT 226.120 105.120 226.410 105.165 ;
        RECT 232.085 105.105 232.405 105.165 ;
        RECT 232.560 105.120 232.850 105.350 ;
        RECT 222.440 104.965 222.730 105.010 ;
        RECT 227.025 104.965 227.345 105.025 ;
        RECT 222.440 104.825 227.345 104.965 ;
        RECT 222.440 104.780 222.730 104.825 ;
        RECT 227.025 104.765 227.345 104.825 ;
        RECT 229.785 104.765 230.105 105.025 ;
        RECT 232.635 104.965 232.775 105.120 ;
        RECT 234.845 105.105 235.165 105.365 ;
        RECT 235.855 105.350 235.995 105.505 ;
        RECT 235.780 105.120 236.070 105.350 ;
        RECT 238.985 105.105 239.305 105.365 ;
        RECT 240.825 105.305 241.145 105.365 ;
        RECT 241.760 105.305 242.050 105.350 ;
        RECT 240.825 105.165 242.050 105.305 ;
        RECT 240.825 105.105 241.145 105.165 ;
        RECT 241.760 105.120 242.050 105.165 ;
        RECT 242.220 105.305 242.510 105.350 ;
        RECT 244.060 105.305 244.350 105.350 ;
        RECT 242.220 105.165 244.350 105.305 ;
        RECT 242.220 105.120 242.510 105.165 ;
        RECT 244.060 105.120 244.350 105.165 ;
        RECT 245.885 105.305 246.205 105.365 ;
        RECT 248.645 105.305 248.965 105.365 ;
        RECT 250.500 105.305 250.790 105.350 ;
        RECT 245.885 105.165 250.790 105.305 ;
        RECT 252.415 105.305 252.555 105.505 ;
        RECT 253.705 105.505 270.035 105.645 ;
        RECT 270.265 105.645 270.585 105.705 ;
        RECT 279.555 105.645 279.695 105.845 ;
        RECT 291.900 105.800 292.190 105.845 ;
        RECT 302.465 105.985 302.785 106.045 ;
        RECT 308.000 105.985 308.290 106.030 ;
        RECT 302.465 105.845 308.290 105.985 ;
        RECT 302.465 105.785 302.785 105.845 ;
        RECT 308.000 105.800 308.290 105.845 ;
        RECT 270.265 105.505 279.695 105.645 ;
        RECT 280.040 105.645 280.330 105.690 ;
        RECT 283.280 105.645 283.930 105.690 ;
        RECT 280.040 105.505 283.930 105.645 ;
        RECT 253.705 105.445 254.025 105.505 ;
        RECT 270.265 105.445 270.585 105.505 ;
        RECT 280.040 105.460 280.630 105.505 ;
        RECT 283.280 105.460 283.930 105.505 ;
        RECT 288.665 105.645 288.985 105.705 ;
        RECT 298.325 105.690 298.645 105.705 ;
        RECT 298.320 105.645 298.970 105.690 ;
        RECT 301.920 105.645 302.210 105.690 ;
        RECT 288.665 105.505 302.210 105.645 ;
        RECT 280.340 105.365 280.630 105.460 ;
        RECT 288.665 105.445 288.985 105.505 ;
        RECT 298.320 105.460 298.970 105.505 ;
        RECT 301.620 105.460 302.210 105.505 ;
        RECT 298.325 105.445 298.645 105.460 ;
        RECT 257.845 105.305 258.165 105.365 ;
        RECT 259.240 105.305 259.530 105.350 ;
        RECT 252.415 105.165 253.475 105.305 ;
        RECT 245.885 105.105 246.205 105.165 ;
        RECT 248.645 105.105 248.965 105.165 ;
        RECT 250.500 105.120 250.790 105.165 ;
        RECT 239.445 104.965 239.765 105.025 ;
        RECT 232.635 104.825 239.765 104.965 ;
        RECT 239.445 104.765 239.765 104.825 ;
        RECT 243.140 104.780 243.430 105.010 ;
        RECT 247.280 104.965 247.570 105.010 ;
        RECT 247.725 104.965 248.045 105.025 ;
        RECT 247.280 104.825 248.045 104.965 ;
        RECT 247.280 104.780 247.570 104.825 ;
        RECT 216.460 104.485 217.135 104.625 ;
        RECT 220.585 104.625 220.905 104.685 ;
        RECT 242.665 104.625 242.985 104.685 ;
        RECT 220.585 104.485 226.335 104.625 ;
        RECT 216.460 104.440 216.750 104.485 ;
        RECT 220.585 104.425 220.905 104.485 ;
        RECT 197.140 104.285 197.430 104.330 ;
        RECT 187.555 104.145 197.430 104.285 ;
        RECT 197.140 104.100 197.430 104.145 ;
        RECT 205.405 104.085 205.725 104.345 ;
        RECT 206.325 104.285 206.645 104.345 ;
        RECT 206.800 104.285 207.090 104.330 ;
        RECT 206.325 104.145 207.090 104.285 ;
        RECT 206.325 104.085 206.645 104.145 ;
        RECT 206.800 104.100 207.090 104.145 ;
        RECT 214.620 104.285 214.910 104.330 ;
        RECT 219.205 104.285 219.525 104.345 ;
        RECT 214.620 104.145 219.525 104.285 ;
        RECT 214.620 104.100 214.910 104.145 ;
        RECT 219.205 104.085 219.525 104.145 ;
        RECT 219.665 104.085 219.985 104.345 ;
        RECT 226.195 104.285 226.335 104.485 ;
        RECT 230.335 104.485 242.985 104.625 ;
        RECT 243.215 104.625 243.355 104.780 ;
        RECT 247.725 104.765 248.045 104.825 ;
        RECT 252.785 104.765 253.105 105.025 ;
        RECT 253.335 104.965 253.475 105.165 ;
        RECT 257.845 105.165 259.530 105.305 ;
        RECT 257.845 105.105 258.165 105.165 ;
        RECT 259.240 105.120 259.530 105.165 ;
        RECT 259.685 105.305 260.005 105.365 ;
        RECT 259.685 105.165 261.295 105.305 ;
        RECT 259.685 105.105 260.005 105.165 ;
        RECT 258.765 104.965 259.085 105.025 ;
        RECT 253.335 104.825 259.085 104.965 ;
        RECT 258.765 104.765 259.085 104.825 ;
        RECT 260.145 104.765 260.465 105.025 ;
        RECT 261.155 104.965 261.295 105.165 ;
        RECT 261.525 105.105 261.845 105.365 ;
        RECT 261.985 105.305 262.305 105.365 ;
        RECT 263.380 105.305 263.670 105.350 ;
        RECT 261.985 105.165 263.670 105.305 ;
        RECT 261.985 105.105 262.305 105.165 ;
        RECT 263.380 105.120 263.670 105.165 ;
        RECT 264.745 105.305 265.065 105.365 ;
        RECT 267.060 105.305 267.350 105.350 ;
        RECT 264.745 105.165 267.350 105.305 ;
        RECT 264.745 105.105 265.065 105.165 ;
        RECT 267.060 105.120 267.350 105.165 ;
        RECT 268.425 105.305 268.745 105.365 ;
        RECT 268.900 105.305 269.190 105.350 ;
        RECT 268.425 105.165 269.190 105.305 ;
        RECT 268.425 105.105 268.745 105.165 ;
        RECT 268.900 105.120 269.190 105.165 ;
        RECT 270.725 105.105 271.045 105.365 ;
        RECT 277.640 105.305 277.930 105.350 ;
        RECT 279.005 105.305 279.325 105.365 ;
        RECT 277.640 105.165 279.325 105.305 ;
        RECT 277.640 105.120 277.930 105.165 ;
        RECT 279.005 105.105 279.325 105.165 ;
        RECT 280.340 105.145 280.705 105.365 ;
        RECT 280.385 105.105 280.705 105.145 ;
        RECT 281.420 105.305 281.710 105.350 ;
        RECT 285.000 105.305 285.290 105.350 ;
        RECT 286.835 105.305 287.125 105.350 ;
        RECT 281.420 105.165 287.125 105.305 ;
        RECT 281.420 105.120 281.710 105.165 ;
        RECT 285.000 105.120 285.290 105.165 ;
        RECT 286.835 105.120 287.125 105.165 ;
        RECT 289.140 105.305 289.430 105.350 ;
        RECT 290.045 105.305 290.365 105.365 ;
        RECT 289.140 105.165 290.365 105.305 ;
        RECT 289.140 105.120 289.430 105.165 ;
        RECT 290.045 105.105 290.365 105.165 ;
        RECT 292.345 105.305 292.665 105.365 ;
        RECT 292.820 105.305 293.110 105.350 ;
        RECT 292.345 105.165 293.110 105.305 ;
        RECT 292.345 105.105 292.665 105.165 ;
        RECT 292.820 105.120 293.110 105.165 ;
        RECT 295.125 105.305 295.415 105.350 ;
        RECT 296.960 105.305 297.250 105.350 ;
        RECT 300.540 105.305 300.830 105.350 ;
        RECT 295.125 105.165 300.830 105.305 ;
        RECT 295.125 105.120 295.415 105.165 ;
        RECT 296.960 105.120 297.250 105.165 ;
        RECT 300.540 105.120 300.830 105.165 ;
        RECT 301.620 105.145 301.910 105.460 ;
        RECT 303.385 105.305 303.705 105.365 ;
        RECT 305.700 105.305 305.990 105.350 ;
        RECT 303.385 105.165 305.990 105.305 ;
        RECT 303.385 105.105 303.705 105.165 ;
        RECT 305.700 105.120 305.990 105.165 ;
        RECT 307.080 105.305 307.370 105.350 ;
        RECT 308.445 105.305 308.765 105.365 ;
        RECT 307.080 105.165 308.765 105.305 ;
        RECT 307.080 105.120 307.370 105.165 ;
        RECT 308.445 105.105 308.765 105.165 ;
        RECT 266.125 104.965 266.445 105.025 ;
        RECT 261.155 104.825 266.445 104.965 ;
        RECT 266.125 104.765 266.445 104.825 ;
        RECT 275.325 104.765 275.645 105.025 ;
        RECT 282.225 104.965 282.545 105.025 ;
        RECT 285.920 104.965 286.210 105.010 ;
        RECT 282.225 104.825 286.210 104.965 ;
        RECT 282.225 104.765 282.545 104.825 ;
        RECT 285.920 104.780 286.210 104.825 ;
        RECT 287.300 104.965 287.590 105.010 ;
        RECT 294.645 104.965 294.965 105.025 ;
        RECT 287.300 104.825 294.965 104.965 ;
        RECT 287.300 104.780 287.590 104.825 ;
        RECT 294.645 104.765 294.965 104.825 ;
        RECT 296.040 104.965 296.330 105.010 ;
        RECT 303.845 104.965 304.165 105.025 ;
        RECT 296.040 104.825 304.165 104.965 ;
        RECT 296.040 104.780 296.330 104.825 ;
        RECT 303.845 104.765 304.165 104.825 ;
        RECT 249.105 104.625 249.425 104.685 ;
        RECT 243.215 104.485 249.425 104.625 ;
        RECT 230.335 104.285 230.475 104.485 ;
        RECT 242.665 104.425 242.985 104.485 ;
        RECT 249.105 104.425 249.425 104.485 ;
        RECT 251.405 104.625 251.725 104.685 ;
        RECT 267.505 104.625 267.825 104.685 ;
        RECT 268.885 104.625 269.205 104.685 ;
        RECT 272.580 104.625 272.870 104.670 ;
        RECT 281.420 104.625 281.710 104.670 ;
        RECT 284.540 104.625 284.830 104.670 ;
        RECT 286.430 104.625 286.720 104.670 ;
        RECT 251.405 104.485 264.975 104.625 ;
        RECT 251.405 104.425 251.725 104.485 ;
        RECT 226.195 104.145 230.475 104.285 ;
        RECT 239.920 104.285 240.210 104.330 ;
        RECT 241.285 104.285 241.605 104.345 ;
        RECT 239.920 104.145 241.605 104.285 ;
        RECT 239.920 104.100 240.210 104.145 ;
        RECT 241.285 104.085 241.605 104.145 ;
        RECT 247.740 104.285 248.030 104.330 ;
        RECT 248.645 104.285 248.965 104.345 ;
        RECT 247.740 104.145 248.965 104.285 ;
        RECT 247.740 104.100 248.030 104.145 ;
        RECT 248.645 104.085 248.965 104.145 ;
        RECT 255.085 104.285 255.405 104.345 ;
        RECT 256.020 104.285 256.310 104.330 ;
        RECT 255.085 104.145 256.310 104.285 ;
        RECT 255.085 104.085 255.405 104.145 ;
        RECT 256.020 104.100 256.310 104.145 ;
        RECT 257.385 104.085 257.705 104.345 ;
        RECT 258.765 104.285 259.085 104.345 ;
        RECT 262.460 104.285 262.750 104.330 ;
        RECT 258.765 104.145 262.750 104.285 ;
        RECT 258.765 104.085 259.085 104.145 ;
        RECT 262.460 104.100 262.750 104.145 ;
        RECT 264.285 104.085 264.605 104.345 ;
        RECT 264.835 104.285 264.975 104.485 ;
        RECT 267.505 104.485 268.655 104.625 ;
        RECT 267.505 104.425 267.825 104.485 ;
        RECT 267.980 104.285 268.270 104.330 ;
        RECT 264.835 104.145 268.270 104.285 ;
        RECT 268.515 104.285 268.655 104.485 ;
        RECT 268.885 104.485 272.870 104.625 ;
        RECT 268.885 104.425 269.205 104.485 ;
        RECT 272.580 104.440 272.870 104.485 ;
        RECT 276.335 104.485 279.235 104.625 ;
        RECT 276.335 104.285 276.475 104.485 ;
        RECT 268.515 104.145 276.475 104.285 ;
        RECT 277.165 104.285 277.485 104.345 ;
        RECT 278.560 104.285 278.850 104.330 ;
        RECT 277.165 104.145 278.850 104.285 ;
        RECT 279.095 104.285 279.235 104.485 ;
        RECT 281.420 104.485 286.720 104.625 ;
        RECT 281.420 104.440 281.710 104.485 ;
        RECT 284.540 104.440 284.830 104.485 ;
        RECT 286.430 104.440 286.720 104.485 ;
        RECT 295.530 104.625 295.820 104.670 ;
        RECT 297.420 104.625 297.710 104.670 ;
        RECT 300.540 104.625 300.830 104.670 ;
        RECT 295.530 104.485 300.830 104.625 ;
        RECT 295.530 104.440 295.820 104.485 ;
        RECT 297.420 104.440 297.710 104.485 ;
        RECT 300.540 104.440 300.830 104.485 ;
        RECT 304.765 104.425 305.085 104.685 ;
        RECT 288.220 104.285 288.510 104.330 ;
        RECT 279.095 104.145 288.510 104.285 ;
        RECT 267.980 104.100 268.270 104.145 ;
        RECT 277.165 104.085 277.485 104.145 ;
        RECT 278.560 104.100 278.850 104.145 ;
        RECT 288.220 104.100 288.510 104.145 ;
        RECT 303.385 104.085 303.705 104.345 ;
        RECT 162.095 103.465 311.135 103.945 ;
        RECT 164.480 103.265 164.770 103.310 ;
        RECT 166.305 103.265 166.625 103.325 ;
        RECT 164.480 103.125 166.625 103.265 ;
        RECT 164.480 103.080 164.770 103.125 ;
        RECT 166.305 103.065 166.625 103.125 ;
        RECT 175.505 103.265 175.825 103.325 ;
        RECT 176.805 103.265 177.095 103.310 ;
        RECT 175.505 103.125 177.095 103.265 ;
        RECT 175.505 103.065 175.825 103.125 ;
        RECT 176.805 103.080 177.095 103.125 ;
        RECT 177.345 103.265 177.665 103.325 ;
        RECT 186.560 103.265 186.850 103.310 ;
        RECT 189.305 103.265 189.625 103.325 ;
        RECT 177.345 103.125 184.475 103.265 ;
        RECT 177.345 103.065 177.665 103.125 ;
        RECT 184.335 102.970 184.475 103.125 ;
        RECT 186.560 103.125 189.625 103.265 ;
        RECT 186.560 103.080 186.850 103.125 ;
        RECT 189.305 103.065 189.625 103.125 ;
        RECT 196.205 103.265 196.525 103.325 ;
        RECT 197.140 103.265 197.430 103.310 ;
        RECT 196.205 103.125 197.430 103.265 ;
        RECT 196.205 103.065 196.525 103.125 ;
        RECT 197.140 103.080 197.430 103.125 ;
        RECT 198.505 103.265 198.825 103.325 ;
        RECT 199.440 103.265 199.730 103.310 ;
        RECT 198.505 103.125 199.730 103.265 ;
        RECT 198.505 103.065 198.825 103.125 ;
        RECT 199.440 103.080 199.730 103.125 ;
        RECT 200.805 103.265 201.125 103.325 ;
        RECT 201.740 103.265 202.030 103.310 ;
        RECT 200.805 103.125 202.030 103.265 ;
        RECT 200.805 103.065 201.125 103.125 ;
        RECT 201.740 103.080 202.030 103.125 ;
        RECT 205.405 103.265 205.725 103.325 ;
        RECT 214.605 103.265 214.925 103.325 ;
        RECT 205.405 103.125 214.925 103.265 ;
        RECT 205.405 103.065 205.725 103.125 ;
        RECT 214.605 103.065 214.925 103.125 ;
        RECT 226.105 103.265 226.425 103.325 ;
        RECT 231.640 103.265 231.930 103.310 ;
        RECT 226.105 103.125 231.930 103.265 ;
        RECT 226.105 103.065 226.425 103.125 ;
        RECT 231.640 103.080 231.930 103.125 ;
        RECT 240.365 103.265 240.685 103.325 ;
        RECT 251.420 103.265 251.710 103.310 ;
        RECT 240.365 103.125 251.710 103.265 ;
        RECT 240.365 103.065 240.685 103.125 ;
        RECT 251.420 103.080 251.710 103.125 ;
        RECT 257.385 103.265 257.705 103.325 ;
        RECT 258.685 103.265 258.975 103.310 ;
        RECT 257.385 103.125 258.975 103.265 ;
        RECT 257.385 103.065 257.705 103.125 ;
        RECT 258.685 103.080 258.975 103.125 ;
        RECT 260.605 103.265 260.925 103.325 ;
        RECT 276.260 103.265 276.550 103.310 ;
        RECT 303.845 103.265 304.165 103.325 ;
        RECT 304.320 103.265 304.610 103.310 ;
        RECT 260.605 103.125 276.550 103.265 ;
        RECT 260.605 103.065 260.925 103.125 ;
        RECT 276.260 103.080 276.550 103.125 ;
        RECT 276.795 103.125 296.255 103.265 ;
        RECT 166.730 102.925 167.020 102.970 ;
        RECT 168.620 102.925 168.910 102.970 ;
        RECT 171.740 102.925 172.030 102.970 ;
        RECT 166.730 102.785 172.030 102.925 ;
        RECT 166.730 102.740 167.020 102.785 ;
        RECT 168.620 102.740 168.910 102.785 ;
        RECT 171.740 102.740 172.030 102.785 ;
        RECT 176.390 102.925 176.680 102.970 ;
        RECT 178.280 102.925 178.570 102.970 ;
        RECT 181.400 102.925 181.690 102.970 ;
        RECT 176.390 102.785 181.690 102.925 ;
        RECT 176.390 102.740 176.680 102.785 ;
        RECT 178.280 102.740 178.570 102.785 ;
        RECT 181.400 102.740 181.690 102.785 ;
        RECT 184.260 102.925 184.550 102.970 ;
        RECT 188.350 102.925 188.640 102.970 ;
        RECT 190.240 102.925 190.530 102.970 ;
        RECT 193.360 102.925 193.650 102.970 ;
        RECT 184.260 102.785 188.155 102.925 ;
        RECT 184.260 102.740 184.550 102.785 ;
        RECT 169.985 102.585 170.305 102.645 ;
        RECT 175.520 102.585 175.810 102.630 ;
        RECT 188.015 102.585 188.155 102.785 ;
        RECT 188.350 102.785 193.650 102.925 ;
        RECT 188.350 102.740 188.640 102.785 ;
        RECT 190.240 102.740 190.530 102.785 ;
        RECT 193.360 102.740 193.650 102.785 ;
        RECT 204.450 102.925 204.740 102.970 ;
        RECT 206.340 102.925 206.630 102.970 ;
        RECT 209.460 102.925 209.750 102.970 ;
        RECT 218.285 102.925 218.605 102.985 ;
        RECT 204.450 102.785 209.750 102.925 ;
        RECT 204.450 102.740 204.740 102.785 ;
        RECT 206.340 102.740 206.630 102.785 ;
        RECT 209.460 102.740 209.750 102.785 ;
        RECT 215.615 102.785 218.605 102.925 ;
        RECT 203.580 102.585 203.870 102.630 ;
        RECT 211.845 102.585 212.165 102.645 ;
        RECT 169.985 102.445 173.205 102.585 ;
        RECT 169.985 102.385 170.305 102.445 ;
        RECT 165.400 102.060 165.690 102.290 ;
        RECT 165.475 101.565 165.615 102.060 ;
        RECT 165.845 102.045 166.165 102.305 ;
        RECT 166.325 102.245 166.615 102.290 ;
        RECT 168.160 102.245 168.450 102.290 ;
        RECT 171.740 102.245 172.030 102.290 ;
        RECT 173.065 102.265 173.205 102.445 ;
        RECT 175.520 102.445 187.695 102.585 ;
        RECT 188.015 102.445 195.515 102.585 ;
        RECT 175.520 102.400 175.810 102.445 ;
        RECT 166.325 102.105 172.030 102.245 ;
        RECT 166.325 102.060 166.615 102.105 ;
        RECT 168.160 102.060 168.450 102.105 ;
        RECT 171.740 102.060 172.030 102.105 ;
        RECT 167.240 101.905 167.530 101.950 ;
        RECT 168.605 101.905 168.925 101.965 ;
        RECT 169.985 101.950 170.305 101.965 ;
        RECT 167.240 101.765 168.925 101.905 ;
        RECT 167.240 101.720 167.530 101.765 ;
        RECT 168.605 101.705 168.925 101.765 ;
        RECT 169.520 101.905 170.305 101.950 ;
        RECT 172.820 101.950 173.205 102.265 ;
        RECT 175.985 102.245 176.275 102.290 ;
        RECT 177.820 102.245 178.110 102.290 ;
        RECT 181.400 102.245 181.690 102.290 ;
        RECT 175.985 102.105 181.690 102.245 ;
        RECT 175.985 102.060 176.275 102.105 ;
        RECT 177.820 102.060 178.110 102.105 ;
        RECT 181.400 102.060 181.690 102.105 ;
        RECT 182.480 101.950 182.770 102.265 ;
        RECT 185.625 102.045 185.945 102.305 ;
        RECT 187.555 102.290 187.695 102.445 ;
        RECT 187.480 102.060 187.770 102.290 ;
        RECT 187.945 102.245 188.235 102.290 ;
        RECT 189.780 102.245 190.070 102.290 ;
        RECT 193.360 102.245 193.650 102.290 ;
        RECT 187.945 102.105 193.650 102.245 ;
        RECT 187.945 102.060 188.235 102.105 ;
        RECT 189.780 102.060 190.070 102.105 ;
        RECT 193.360 102.060 193.650 102.105 ;
        RECT 172.820 101.905 173.410 101.950 ;
        RECT 179.180 101.905 179.830 101.950 ;
        RECT 182.480 101.905 183.070 101.950 ;
        RECT 187.555 101.905 187.695 102.060 ;
        RECT 188.385 101.905 188.705 101.965 ;
        RECT 169.520 101.765 183.070 101.905 ;
        RECT 169.520 101.720 170.305 101.765 ;
        RECT 173.120 101.720 173.410 101.765 ;
        RECT 169.985 101.705 170.305 101.720 ;
        RECT 174.125 101.565 174.445 101.625 ;
        RECT 165.475 101.425 174.445 101.565 ;
        RECT 174.125 101.365 174.445 101.425 ;
        RECT 174.585 101.565 174.905 101.625 ;
        RECT 176.885 101.565 177.205 101.625 ;
        RECT 174.585 101.425 177.205 101.565 ;
        RECT 178.815 101.565 178.955 101.765 ;
        RECT 179.180 101.720 179.830 101.765 ;
        RECT 182.780 101.720 183.070 101.765 ;
        RECT 183.875 101.765 187.235 101.905 ;
        RECT 187.555 101.765 188.705 101.905 ;
        RECT 183.875 101.565 184.015 101.765 ;
        RECT 178.815 101.425 184.015 101.565 ;
        RECT 187.095 101.565 187.235 101.765 ;
        RECT 188.385 101.705 188.705 101.765 ;
        RECT 188.845 101.705 189.165 101.965 ;
        RECT 191.145 101.950 191.465 101.965 ;
        RECT 194.440 101.950 194.730 102.265 ;
        RECT 191.140 101.905 191.790 101.950 ;
        RECT 194.440 101.905 195.030 101.950 ;
        RECT 189.395 101.765 195.030 101.905 ;
        RECT 195.375 101.905 195.515 102.445 ;
        RECT 203.580 102.445 212.165 102.585 ;
        RECT 203.580 102.400 203.870 102.445 ;
        RECT 211.845 102.385 212.165 102.445 ;
        RECT 212.320 102.585 212.610 102.630 ;
        RECT 212.765 102.585 213.085 102.645 ;
        RECT 215.615 102.630 215.755 102.785 ;
        RECT 218.285 102.725 218.605 102.785 ;
        RECT 220.240 102.925 220.530 102.970 ;
        RECT 223.360 102.925 223.650 102.970 ;
        RECT 225.250 102.925 225.540 102.970 ;
        RECT 227.040 102.925 227.330 102.970 ;
        RECT 220.240 102.785 225.540 102.925 ;
        RECT 220.240 102.740 220.530 102.785 ;
        RECT 223.360 102.740 223.650 102.785 ;
        RECT 225.250 102.740 225.540 102.785 ;
        RECT 226.195 102.785 227.330 102.925 ;
        RECT 212.320 102.445 213.085 102.585 ;
        RECT 212.320 102.400 212.610 102.445 ;
        RECT 212.765 102.385 213.085 102.445 ;
        RECT 215.540 102.400 215.830 102.630 ;
        RECT 221.965 102.585 222.285 102.645 ;
        RECT 216.075 102.445 222.285 102.585 ;
        RECT 197.585 102.245 197.905 102.305 ;
        RECT 198.060 102.245 198.350 102.290 ;
        RECT 197.585 102.105 198.350 102.245 ;
        RECT 197.585 102.045 197.905 102.105 ;
        RECT 198.060 102.060 198.350 102.105 ;
        RECT 199.425 102.245 199.745 102.305 ;
        RECT 200.360 102.245 200.650 102.290 ;
        RECT 199.425 102.105 200.650 102.245 ;
        RECT 199.425 102.045 199.745 102.105 ;
        RECT 200.360 102.060 200.650 102.105 ;
        RECT 202.645 102.045 202.965 102.305 ;
        RECT 204.045 102.245 204.335 102.290 ;
        RECT 205.880 102.245 206.170 102.290 ;
        RECT 209.460 102.245 209.750 102.290 ;
        RECT 204.045 102.105 209.750 102.245 ;
        RECT 204.045 102.060 204.335 102.105 ;
        RECT 205.880 102.060 206.170 102.105 ;
        RECT 209.460 102.060 209.750 102.105 ;
        RECT 210.005 102.245 210.325 102.305 ;
        RECT 210.540 102.245 210.830 102.265 ;
        RECT 216.075 102.245 216.215 102.445 ;
        RECT 221.965 102.385 222.285 102.445 ;
        RECT 224.740 102.585 225.030 102.630 ;
        RECT 226.195 102.585 226.335 102.785 ;
        RECT 227.040 102.740 227.330 102.785 ;
        RECT 238.030 102.925 238.320 102.970 ;
        RECT 239.920 102.925 240.210 102.970 ;
        RECT 243.040 102.925 243.330 102.970 ;
        RECT 238.030 102.785 243.330 102.925 ;
        RECT 238.030 102.740 238.320 102.785 ;
        RECT 239.920 102.740 240.210 102.785 ;
        RECT 243.040 102.740 243.330 102.785 ;
        RECT 245.885 102.725 246.205 102.985 ;
        RECT 246.360 102.740 246.650 102.970 ;
        RECT 258.270 102.925 258.560 102.970 ;
        RECT 260.160 102.925 260.450 102.970 ;
        RECT 263.280 102.925 263.570 102.970 ;
        RECT 249.195 102.785 255.775 102.925 ;
        RECT 224.740 102.445 226.335 102.585 ;
        RECT 227.485 102.585 227.805 102.645 ;
        RECT 229.800 102.585 230.090 102.630 ;
        RECT 237.160 102.585 237.450 102.630 ;
        RECT 227.485 102.445 230.090 102.585 ;
        RECT 224.740 102.400 225.030 102.445 ;
        RECT 227.485 102.385 227.805 102.445 ;
        RECT 229.800 102.400 230.090 102.445 ;
        RECT 230.335 102.445 237.450 102.585 ;
        RECT 210.005 102.105 216.215 102.245 ;
        RECT 210.005 102.045 210.325 102.105 ;
        RECT 203.565 101.905 203.885 101.965 ;
        RECT 195.375 101.765 203.885 101.905 ;
        RECT 189.395 101.565 189.535 101.765 ;
        RECT 191.140 101.720 191.790 101.765 ;
        RECT 194.740 101.720 195.030 101.765 ;
        RECT 191.145 101.705 191.465 101.720 ;
        RECT 203.565 101.705 203.885 101.765 ;
        RECT 204.960 101.905 205.250 101.950 ;
        RECT 206.325 101.905 206.645 101.965 ;
        RECT 210.540 101.950 210.830 102.105 ;
        RECT 219.160 101.950 219.450 102.265 ;
        RECT 220.240 102.245 220.530 102.290 ;
        RECT 223.820 102.245 224.110 102.290 ;
        RECT 225.655 102.245 225.945 102.290 ;
        RECT 220.240 102.105 225.945 102.245 ;
        RECT 220.240 102.060 220.530 102.105 ;
        RECT 223.820 102.060 224.110 102.105 ;
        RECT 225.655 102.060 225.945 102.105 ;
        RECT 226.105 102.245 226.425 102.305 ;
        RECT 230.335 102.245 230.475 102.445 ;
        RECT 237.160 102.400 237.450 102.445 ;
        RECT 238.540 102.585 238.830 102.630 ;
        RECT 246.435 102.585 246.575 102.740 ;
        RECT 249.195 102.645 249.335 102.785 ;
        RECT 238.540 102.445 246.575 102.585 ;
        RECT 238.540 102.400 238.830 102.445 ;
        RECT 248.645 102.385 248.965 102.645 ;
        RECT 249.105 102.385 249.425 102.645 ;
        RECT 255.085 102.385 255.405 102.645 ;
        RECT 255.635 102.630 255.775 102.785 ;
        RECT 258.270 102.785 263.570 102.925 ;
        RECT 258.270 102.740 258.560 102.785 ;
        RECT 260.160 102.740 260.450 102.785 ;
        RECT 263.280 102.740 263.570 102.785 ;
        RECT 266.125 102.725 266.445 102.985 ;
        RECT 267.470 102.925 267.760 102.970 ;
        RECT 269.360 102.925 269.650 102.970 ;
        RECT 272.480 102.925 272.770 102.970 ;
        RECT 267.470 102.785 272.770 102.925 ;
        RECT 267.470 102.740 267.760 102.785 ;
        RECT 269.360 102.740 269.650 102.785 ;
        RECT 272.480 102.740 272.770 102.785 ;
        RECT 255.560 102.400 255.850 102.630 ;
        RECT 266.600 102.585 266.890 102.630 ;
        RECT 269.805 102.585 270.125 102.645 ;
        RECT 257.475 102.445 270.125 102.585 ;
        RECT 226.105 102.105 230.475 102.245 ;
        RECT 226.105 102.045 226.425 102.105 ;
        RECT 232.545 102.045 232.865 102.305 ;
        RECT 237.625 102.245 237.915 102.290 ;
        RECT 239.460 102.245 239.750 102.290 ;
        RECT 243.040 102.245 243.330 102.290 ;
        RECT 237.625 102.105 243.330 102.245 ;
        RECT 237.625 102.060 237.915 102.105 ;
        RECT 239.460 102.060 239.750 102.105 ;
        RECT 243.040 102.060 243.330 102.105 ;
        RECT 204.960 101.765 206.645 101.905 ;
        RECT 204.960 101.720 205.250 101.765 ;
        RECT 206.325 101.705 206.645 101.765 ;
        RECT 207.240 101.905 207.890 101.950 ;
        RECT 210.540 101.905 211.130 101.950 ;
        RECT 207.240 101.765 211.130 101.905 ;
        RECT 207.240 101.720 207.890 101.765 ;
        RECT 210.840 101.720 211.130 101.765 ;
        RECT 218.860 101.905 219.450 101.950 ;
        RECT 221.965 101.950 222.285 101.965 ;
        RECT 221.965 101.905 222.750 101.950 ;
        RECT 218.860 101.765 222.750 101.905 ;
        RECT 218.860 101.720 219.150 101.765 ;
        RECT 221.965 101.720 222.750 101.765 ;
        RECT 228.405 101.905 228.725 101.965 ;
        RECT 229.325 101.905 229.645 101.965 ;
        RECT 244.120 101.950 244.410 102.265 ;
        RECT 247.725 102.245 248.045 102.305 ;
        RECT 250.500 102.245 250.790 102.290 ;
        RECT 247.725 102.105 250.790 102.245 ;
        RECT 247.725 102.045 248.045 102.105 ;
        RECT 250.500 102.060 250.790 102.105 ;
        RECT 254.625 102.045 254.945 102.305 ;
        RECT 255.635 102.245 255.775 102.400 ;
        RECT 257.475 102.305 257.615 102.445 ;
        RECT 266.600 102.400 266.890 102.445 ;
        RECT 269.805 102.385 270.125 102.445 ;
        RECT 255.635 102.105 257.155 102.245 ;
        RECT 228.405 101.765 229.645 101.905 ;
        RECT 221.965 101.705 222.285 101.720 ;
        RECT 228.405 101.705 228.725 101.765 ;
        RECT 229.325 101.705 229.645 101.765 ;
        RECT 240.820 101.905 241.470 101.950 ;
        RECT 244.120 101.905 244.710 101.950 ;
        RECT 246.345 101.905 246.665 101.965 ;
        RECT 257.015 101.905 257.155 102.105 ;
        RECT 257.385 102.045 257.705 102.305 ;
        RECT 257.865 102.245 258.155 102.290 ;
        RECT 259.700 102.245 259.990 102.290 ;
        RECT 263.280 102.245 263.570 102.290 ;
        RECT 257.865 102.105 263.570 102.245 ;
        RECT 257.865 102.060 258.155 102.105 ;
        RECT 259.700 102.060 259.990 102.105 ;
        RECT 263.280 102.060 263.570 102.105 ;
        RECT 260.145 101.905 260.465 101.965 ;
        RECT 264.360 101.950 264.650 102.265 ;
        RECT 267.065 102.245 267.355 102.290 ;
        RECT 268.900 102.245 269.190 102.290 ;
        RECT 272.480 102.245 272.770 102.290 ;
        RECT 267.065 102.105 272.770 102.245 ;
        RECT 267.065 102.060 267.355 102.105 ;
        RECT 268.900 102.060 269.190 102.105 ;
        RECT 272.480 102.060 272.770 102.105 ;
        RECT 273.560 102.245 273.850 102.265 ;
        RECT 276.795 102.245 276.935 103.125 ;
        RECT 281.420 102.925 281.710 102.970 ;
        RECT 284.540 102.925 284.830 102.970 ;
        RECT 286.430 102.925 286.720 102.970 ;
        RECT 288.665 102.925 288.985 102.985 ;
        RECT 281.420 102.785 286.720 102.925 ;
        RECT 281.420 102.740 281.710 102.785 ;
        RECT 284.540 102.740 284.830 102.785 ;
        RECT 286.430 102.740 286.720 102.785 ;
        RECT 286.915 102.785 288.985 102.925 ;
        RECT 286.915 102.585 287.055 102.785 ;
        RECT 288.665 102.725 288.985 102.785 ;
        RECT 290.620 102.925 290.910 102.970 ;
        RECT 293.740 102.925 294.030 102.970 ;
        RECT 295.630 102.925 295.920 102.970 ;
        RECT 290.620 102.785 295.920 102.925 ;
        RECT 296.115 102.925 296.255 103.125 ;
        RECT 303.845 103.125 304.610 103.265 ;
        RECT 303.845 103.065 304.165 103.125 ;
        RECT 304.320 103.080 304.610 103.125 ;
        RECT 305.225 102.925 305.545 102.985 ;
        RECT 296.115 102.785 305.545 102.925 ;
        RECT 290.620 102.740 290.910 102.785 ;
        RECT 293.740 102.740 294.030 102.785 ;
        RECT 295.630 102.740 295.920 102.785 ;
        RECT 305.225 102.725 305.545 102.785 ;
        RECT 294.645 102.585 294.965 102.645 ;
        RECT 280.475 102.445 287.055 102.585 ;
        RECT 287.835 102.445 294.965 102.585 ;
        RECT 280.475 102.305 280.615 102.445 ;
        RECT 273.560 102.105 276.935 102.245 ;
        RECT 240.820 101.765 253.475 101.905 ;
        RECT 257.015 101.765 260.465 101.905 ;
        RECT 240.820 101.720 241.470 101.765 ;
        RECT 244.420 101.720 244.710 101.765 ;
        RECT 246.345 101.705 246.665 101.765 ;
        RECT 187.095 101.425 189.535 101.565 ;
        RECT 174.585 101.365 174.905 101.425 ;
        RECT 176.885 101.365 177.205 101.425 ;
        RECT 196.205 101.365 196.525 101.625 ;
        RECT 212.765 101.365 213.085 101.625 ;
        RECT 213.685 101.565 214.005 101.625 ;
        RECT 214.620 101.565 214.910 101.610 ;
        RECT 213.685 101.425 214.910 101.565 ;
        RECT 213.685 101.365 214.005 101.425 ;
        RECT 214.620 101.380 214.910 101.425 ;
        RECT 215.065 101.365 215.385 101.625 ;
        RECT 217.365 101.365 217.685 101.625 ;
        RECT 228.880 101.565 229.170 101.610 ;
        RECT 229.785 101.565 230.105 101.625 ;
        RECT 228.880 101.425 230.105 101.565 ;
        RECT 228.880 101.380 229.170 101.425 ;
        RECT 229.785 101.365 230.105 101.425 ;
        RECT 242.665 101.565 242.985 101.625 ;
        RECT 248.185 101.565 248.505 101.625 ;
        RECT 242.665 101.425 248.505 101.565 ;
        RECT 242.665 101.365 242.985 101.425 ;
        RECT 248.185 101.365 248.505 101.425 ;
        RECT 251.865 101.565 252.185 101.625 ;
        RECT 252.800 101.565 253.090 101.610 ;
        RECT 251.865 101.425 253.090 101.565 ;
        RECT 253.335 101.565 253.475 101.765 ;
        RECT 260.145 101.705 260.465 101.765 ;
        RECT 261.060 101.905 261.710 101.950 ;
        RECT 264.360 101.905 264.950 101.950 ;
        RECT 261.060 101.765 265.435 101.905 ;
        RECT 261.060 101.720 261.710 101.765 ;
        RECT 264.660 101.720 264.950 101.765 ;
        RECT 257.845 101.565 258.165 101.625 ;
        RECT 265.295 101.565 265.435 101.765 ;
        RECT 267.965 101.705 268.285 101.965 ;
        RECT 273.560 101.950 273.850 102.105 ;
        RECT 277.165 102.045 277.485 102.305 ;
        RECT 280.385 102.265 280.705 102.305 ;
        RECT 280.340 102.045 280.705 102.265 ;
        RECT 281.420 102.245 281.710 102.290 ;
        RECT 285.000 102.245 285.290 102.290 ;
        RECT 286.835 102.245 287.125 102.290 ;
        RECT 281.420 102.105 287.125 102.245 ;
        RECT 281.420 102.060 281.710 102.105 ;
        RECT 285.000 102.060 285.290 102.105 ;
        RECT 286.835 102.060 287.125 102.105 ;
        RECT 287.300 102.245 287.590 102.290 ;
        RECT 287.835 102.245 287.975 102.445 ;
        RECT 294.645 102.385 294.965 102.445 ;
        RECT 295.105 102.585 295.425 102.645 ;
        RECT 296.500 102.585 296.790 102.630 ;
        RECT 295.105 102.445 296.790 102.585 ;
        RECT 295.105 102.385 295.425 102.445 ;
        RECT 296.500 102.400 296.790 102.445 ;
        RECT 297.865 102.585 298.185 102.645 ;
        RECT 299.720 102.585 300.010 102.630 ;
        RECT 307.080 102.585 307.370 102.630 ;
        RECT 297.865 102.445 307.370 102.585 ;
        RECT 297.865 102.385 298.185 102.445 ;
        RECT 299.720 102.400 300.010 102.445 ;
        RECT 307.080 102.400 307.370 102.445 ;
        RECT 287.300 102.105 287.975 102.245 ;
        RECT 287.300 102.060 287.590 102.105 ;
        RECT 270.260 101.905 270.910 101.950 ;
        RECT 273.560 101.905 274.150 101.950 ;
        RECT 270.260 101.765 274.150 101.905 ;
        RECT 270.260 101.720 270.910 101.765 ;
        RECT 273.575 101.565 273.715 101.765 ;
        RECT 273.860 101.720 274.150 101.765 ;
        RECT 274.405 101.905 274.725 101.965 ;
        RECT 280.340 101.950 280.630 102.045 ;
        RECT 280.040 101.905 280.630 101.950 ;
        RECT 283.280 101.905 283.930 101.950 ;
        RECT 274.405 101.765 279.695 101.905 ;
        RECT 274.405 101.705 274.725 101.765 ;
        RECT 253.335 101.425 273.715 101.565 ;
        RECT 251.865 101.365 252.185 101.425 ;
        RECT 252.800 101.380 253.090 101.425 ;
        RECT 257.845 101.365 258.165 101.425 ;
        RECT 275.325 101.365 275.645 101.625 ;
        RECT 277.625 101.565 277.945 101.625 ;
        RECT 278.560 101.565 278.850 101.610 ;
        RECT 277.625 101.425 278.850 101.565 ;
        RECT 279.555 101.565 279.695 101.765 ;
        RECT 280.040 101.765 283.930 101.905 ;
        RECT 280.040 101.720 280.330 101.765 ;
        RECT 283.280 101.720 283.930 101.765 ;
        RECT 285.905 101.705 286.225 101.965 ;
        RECT 288.665 101.905 288.985 101.965 ;
        RECT 289.540 101.950 289.830 102.265 ;
        RECT 290.620 102.245 290.910 102.290 ;
        RECT 294.200 102.245 294.490 102.290 ;
        RECT 296.035 102.245 296.325 102.290 ;
        RECT 290.620 102.105 296.325 102.245 ;
        RECT 290.620 102.060 290.910 102.105 ;
        RECT 294.200 102.060 294.490 102.105 ;
        RECT 296.035 102.060 296.325 102.105 ;
        RECT 302.465 102.045 302.785 102.305 ;
        RECT 303.385 102.245 303.705 102.305 ;
        RECT 306.160 102.245 306.450 102.290 ;
        RECT 303.385 102.105 306.450 102.245 ;
        RECT 303.385 102.045 303.705 102.105 ;
        RECT 306.160 102.060 306.450 102.105 ;
        RECT 289.240 101.905 289.830 101.950 ;
        RECT 292.480 101.905 293.130 101.950 ;
        RECT 287.375 101.765 288.435 101.905 ;
        RECT 287.375 101.565 287.515 101.765 ;
        RECT 279.555 101.425 287.515 101.565 ;
        RECT 277.625 101.365 277.945 101.425 ;
        RECT 278.560 101.380 278.850 101.425 ;
        RECT 287.745 101.365 288.065 101.625 ;
        RECT 288.295 101.565 288.435 101.765 ;
        RECT 288.665 101.765 293.130 101.905 ;
        RECT 288.665 101.705 288.985 101.765 ;
        RECT 289.240 101.720 289.530 101.765 ;
        RECT 292.480 101.720 293.130 101.765 ;
        RECT 293.725 101.905 294.045 101.965 ;
        RECT 295.120 101.905 295.410 101.950 ;
        RECT 293.725 101.765 295.410 101.905 ;
        RECT 293.725 101.705 294.045 101.765 ;
        RECT 295.120 101.720 295.410 101.765 ;
        RECT 295.655 101.765 301.775 101.905 ;
        RECT 295.655 101.565 295.795 101.765 ;
        RECT 288.295 101.425 295.795 101.565 ;
        RECT 296.485 101.565 296.805 101.625 ;
        RECT 296.960 101.565 297.250 101.610 ;
        RECT 296.485 101.425 297.250 101.565 ;
        RECT 296.485 101.365 296.805 101.425 ;
        RECT 296.960 101.380 297.250 101.425 ;
        RECT 298.325 101.565 298.645 101.625 ;
        RECT 298.800 101.565 299.090 101.610 ;
        RECT 298.325 101.425 299.090 101.565 ;
        RECT 298.325 101.365 298.645 101.425 ;
        RECT 298.800 101.380 299.090 101.425 ;
        RECT 299.245 101.365 299.565 101.625 ;
        RECT 301.635 101.610 301.775 101.765 ;
        RECT 301.560 101.380 301.850 101.610 ;
        RECT 306.620 101.565 306.910 101.610 ;
        RECT 307.065 101.565 307.385 101.625 ;
        RECT 306.620 101.425 307.385 101.565 ;
        RECT 306.620 101.380 306.910 101.425 ;
        RECT 307.065 101.365 307.385 101.425 ;
        RECT 162.095 100.745 311.135 101.225 ;
        RECT 164.005 100.545 164.325 100.605 ;
        RECT 164.940 100.545 165.230 100.590 ;
        RECT 164.005 100.405 165.230 100.545 ;
        RECT 164.005 100.345 164.325 100.405 ;
        RECT 164.940 100.360 165.230 100.405 ;
        RECT 175.980 100.545 176.270 100.590 ;
        RECT 182.420 100.545 182.710 100.590 ;
        RECT 182.865 100.545 183.185 100.605 ;
        RECT 175.980 100.405 178.955 100.545 ;
        RECT 175.980 100.360 176.270 100.405 ;
        RECT 169.985 100.205 170.305 100.265 ;
        RECT 170.900 100.205 171.550 100.250 ;
        RECT 174.500 100.205 174.790 100.250 ;
        RECT 169.985 100.065 174.790 100.205 ;
        RECT 169.985 100.005 170.305 100.065 ;
        RECT 170.900 100.020 171.550 100.065 ;
        RECT 174.200 100.020 174.790 100.065 ;
        RECT 165.860 99.865 166.150 99.910 ;
        RECT 166.305 99.865 166.625 99.925 ;
        RECT 165.860 99.725 166.625 99.865 ;
        RECT 165.860 99.680 166.150 99.725 ;
        RECT 166.305 99.665 166.625 99.725 ;
        RECT 167.705 99.865 167.995 99.910 ;
        RECT 169.540 99.865 169.830 99.910 ;
        RECT 173.120 99.865 173.410 99.910 ;
        RECT 167.705 99.725 173.410 99.865 ;
        RECT 167.705 99.680 167.995 99.725 ;
        RECT 169.540 99.680 169.830 99.725 ;
        RECT 173.120 99.680 173.410 99.725 ;
        RECT 174.200 99.705 174.490 100.020 ;
        RECT 178.815 99.910 178.955 100.405 ;
        RECT 182.420 100.405 183.185 100.545 ;
        RECT 182.420 100.360 182.710 100.405 ;
        RECT 182.865 100.345 183.185 100.405 ;
        RECT 184.245 100.545 184.565 100.605 ;
        RECT 185.640 100.545 185.930 100.590 ;
        RECT 184.245 100.405 185.930 100.545 ;
        RECT 184.245 100.345 184.565 100.405 ;
        RECT 185.640 100.360 185.930 100.405 ;
        RECT 187.480 100.545 187.770 100.590 ;
        RECT 189.765 100.545 190.085 100.605 ;
        RECT 187.480 100.405 190.085 100.545 ;
        RECT 187.480 100.360 187.770 100.405 ;
        RECT 189.765 100.345 190.085 100.405 ;
        RECT 197.140 100.545 197.430 100.590 ;
        RECT 198.965 100.545 199.285 100.605 ;
        RECT 197.140 100.405 199.655 100.545 ;
        RECT 197.140 100.360 197.430 100.405 ;
        RECT 198.965 100.345 199.285 100.405 ;
        RECT 179.200 100.205 179.490 100.250 ;
        RECT 185.165 100.205 185.485 100.265 ;
        RECT 190.225 100.205 190.545 100.265 ;
        RECT 179.200 100.065 190.545 100.205 ;
        RECT 179.200 100.020 179.490 100.065 ;
        RECT 185.165 100.005 185.485 100.065 ;
        RECT 190.225 100.005 190.545 100.065 ;
        RECT 191.145 100.205 191.465 100.265 ;
        RECT 192.060 100.205 192.710 100.250 ;
        RECT 195.660 100.205 195.950 100.250 ;
        RECT 191.145 100.065 195.950 100.205 ;
        RECT 191.145 100.005 191.465 100.065 ;
        RECT 192.060 100.020 192.710 100.065 ;
        RECT 195.360 100.020 195.950 100.065 ;
        RECT 178.740 99.865 179.030 99.910 ;
        RECT 183.340 99.865 183.630 99.910 ;
        RECT 183.785 99.865 184.105 99.925 ;
        RECT 178.740 99.725 184.105 99.865 ;
        RECT 178.740 99.680 179.030 99.725 ;
        RECT 183.340 99.680 183.630 99.725 ;
        RECT 183.785 99.665 184.105 99.725 ;
        RECT 188.865 99.865 189.155 99.910 ;
        RECT 190.700 99.865 190.990 99.910 ;
        RECT 194.280 99.865 194.570 99.910 ;
        RECT 188.865 99.725 194.570 99.865 ;
        RECT 188.865 99.680 189.155 99.725 ;
        RECT 190.700 99.680 190.990 99.725 ;
        RECT 194.280 99.680 194.570 99.725 ;
        RECT 195.360 99.705 195.650 100.020 ;
        RECT 199.515 99.910 199.655 100.405 ;
        RECT 199.885 100.345 200.205 100.605 ;
        RECT 212.305 100.545 212.625 100.605 ;
        RECT 214.620 100.545 214.910 100.590 ;
        RECT 212.305 100.405 214.910 100.545 ;
        RECT 212.305 100.345 212.625 100.405 ;
        RECT 214.620 100.360 214.910 100.405 ;
        RECT 226.565 100.345 226.885 100.605 ;
        RECT 227.025 100.345 227.345 100.605 ;
        RECT 257.385 100.545 257.705 100.605 ;
        RECT 239.995 100.405 257.705 100.545 ;
        RECT 204.600 100.205 204.890 100.250 ;
        RECT 207.840 100.205 208.490 100.250 ;
        RECT 210.005 100.205 210.325 100.265 ;
        RECT 204.600 100.065 210.325 100.205 ;
        RECT 204.600 100.020 205.190 100.065 ;
        RECT 207.840 100.020 208.490 100.065 ;
        RECT 199.440 99.865 199.730 99.910 ;
        RECT 199.440 99.725 203.795 99.865 ;
        RECT 199.440 99.680 199.730 99.725 ;
        RECT 167.225 99.325 167.545 99.585 ;
        RECT 168.620 99.525 168.910 99.570 ;
        RECT 168.620 99.385 177.115 99.525 ;
        RECT 168.620 99.340 168.910 99.385 ;
        RECT 176.975 99.230 177.115 99.385 ;
        RECT 179.645 99.325 179.965 99.585 ;
        RECT 184.720 99.340 185.010 99.570 ;
        RECT 185.180 99.525 185.470 99.570 ;
        RECT 186.085 99.525 186.405 99.585 ;
        RECT 185.180 99.385 186.405 99.525 ;
        RECT 185.180 99.340 185.470 99.385 ;
        RECT 168.110 99.185 168.400 99.230 ;
        RECT 170.000 99.185 170.290 99.230 ;
        RECT 173.120 99.185 173.410 99.230 ;
        RECT 168.110 99.045 173.410 99.185 ;
        RECT 168.110 99.000 168.400 99.045 ;
        RECT 170.000 99.000 170.290 99.045 ;
        RECT 173.120 99.000 173.410 99.045 ;
        RECT 176.900 99.000 177.190 99.230 ;
        RECT 184.795 99.185 184.935 99.340 ;
        RECT 186.085 99.325 186.405 99.385 ;
        RECT 188.385 99.325 188.705 99.585 ;
        RECT 189.780 99.525 190.070 99.570 ;
        RECT 189.780 99.385 197.815 99.525 ;
        RECT 189.780 99.340 190.070 99.385 ;
        RECT 197.675 99.230 197.815 99.385 ;
        RECT 200.345 99.325 200.665 99.585 ;
        RECT 203.655 99.525 203.795 99.725 ;
        RECT 204.900 99.705 205.190 100.020 ;
        RECT 210.005 100.005 210.325 100.065 ;
        RECT 210.480 100.205 210.770 100.250 ;
        RECT 212.765 100.205 213.085 100.265 ;
        RECT 210.480 100.065 213.085 100.205 ;
        RECT 210.480 100.020 210.770 100.065 ;
        RECT 212.765 100.005 213.085 100.065 ;
        RECT 219.220 100.205 219.510 100.250 ;
        RECT 219.665 100.205 219.985 100.265 ;
        RECT 221.965 100.250 222.285 100.265 ;
        RECT 219.220 100.065 219.985 100.205 ;
        RECT 219.220 100.020 219.510 100.065 ;
        RECT 219.665 100.005 219.985 100.065 ;
        RECT 221.500 100.205 222.285 100.250 ;
        RECT 225.100 100.205 225.390 100.250 ;
        RECT 221.500 100.065 225.390 100.205 ;
        RECT 226.655 100.205 226.795 100.345 ;
        RECT 228.865 100.205 229.185 100.265 ;
        RECT 226.655 100.065 229.185 100.205 ;
        RECT 221.500 100.020 222.285 100.065 ;
        RECT 221.965 100.005 222.285 100.020 ;
        RECT 224.800 100.020 225.390 100.065 ;
        RECT 205.980 99.865 206.270 99.910 ;
        RECT 209.560 99.865 209.850 99.910 ;
        RECT 211.395 99.865 211.685 99.910 ;
        RECT 205.980 99.725 211.685 99.865 ;
        RECT 205.980 99.680 206.270 99.725 ;
        RECT 209.560 99.680 209.850 99.725 ;
        RECT 211.395 99.680 211.685 99.725 ;
        RECT 215.525 99.665 215.845 99.925 ;
        RECT 218.305 99.865 218.595 99.910 ;
        RECT 220.140 99.865 220.430 99.910 ;
        RECT 223.720 99.865 224.010 99.910 ;
        RECT 218.305 99.725 224.010 99.865 ;
        RECT 218.305 99.680 218.595 99.725 ;
        RECT 220.140 99.680 220.430 99.725 ;
        RECT 223.720 99.680 224.010 99.725 ;
        RECT 224.800 99.705 225.090 100.020 ;
        RECT 228.865 100.005 229.185 100.065 ;
        RECT 227.945 99.665 228.265 99.925 ;
        RECT 239.995 99.910 240.135 100.405 ;
        RECT 241.285 100.005 241.605 100.265 ;
        RECT 243.580 100.205 244.230 100.250 ;
        RECT 246.345 100.205 246.665 100.265 ;
        RECT 247.180 100.205 247.470 100.250 ;
        RECT 243.580 100.065 247.470 100.205 ;
        RECT 243.580 100.020 244.230 100.065 ;
        RECT 246.345 100.005 246.665 100.065 ;
        RECT 246.880 100.020 247.470 100.065 ;
        RECT 239.920 99.680 240.210 99.910 ;
        RECT 240.385 99.865 240.675 99.910 ;
        RECT 242.220 99.865 242.510 99.910 ;
        RECT 245.800 99.865 246.090 99.910 ;
        RECT 240.385 99.725 246.090 99.865 ;
        RECT 240.385 99.680 240.675 99.725 ;
        RECT 242.220 99.680 242.510 99.725 ;
        RECT 245.800 99.680 246.090 99.725 ;
        RECT 246.880 99.705 247.170 100.020 ;
        RECT 249.195 99.910 249.335 100.405 ;
        RECT 257.385 100.345 257.705 100.405 ;
        RECT 258.780 100.360 259.070 100.590 ;
        RECT 267.060 100.545 267.350 100.590 ;
        RECT 267.965 100.545 268.285 100.605 ;
        RECT 267.060 100.405 268.285 100.545 ;
        RECT 267.060 100.360 267.350 100.405 ;
        RECT 250.500 100.205 250.790 100.250 ;
        RECT 251.865 100.205 252.185 100.265 ;
        RECT 250.500 100.065 252.185 100.205 ;
        RECT 250.500 100.020 250.790 100.065 ;
        RECT 251.865 100.005 252.185 100.065 ;
        RECT 252.780 100.205 253.430 100.250 ;
        RECT 256.380 100.205 256.670 100.250 ;
        RECT 257.845 100.205 258.165 100.265 ;
        RECT 252.780 100.065 258.165 100.205 ;
        RECT 252.780 100.020 253.430 100.065 ;
        RECT 256.080 100.020 256.670 100.065 ;
        RECT 249.120 99.680 249.410 99.910 ;
        RECT 249.585 99.865 249.875 99.910 ;
        RECT 251.420 99.865 251.710 99.910 ;
        RECT 255.000 99.865 255.290 99.910 ;
        RECT 249.585 99.725 255.290 99.865 ;
        RECT 249.585 99.680 249.875 99.725 ;
        RECT 251.420 99.680 251.710 99.725 ;
        RECT 255.000 99.680 255.290 99.725 ;
        RECT 256.080 99.705 256.370 100.020 ;
        RECT 257.845 100.005 258.165 100.065 ;
        RECT 258.855 99.865 258.995 100.360 ;
        RECT 267.965 100.345 268.285 100.405 ;
        RECT 268.885 100.345 269.205 100.605 ;
        RECT 277.625 100.545 277.945 100.605 ;
        RECT 281.765 100.545 282.085 100.605 ;
        RECT 282.700 100.545 282.990 100.590 ;
        RECT 277.625 100.405 282.990 100.545 ;
        RECT 277.625 100.345 277.945 100.405 ;
        RECT 281.765 100.345 282.085 100.405 ;
        RECT 282.700 100.360 282.990 100.405 ;
        RECT 284.540 100.545 284.830 100.590 ;
        RECT 285.905 100.545 286.225 100.605 ;
        RECT 284.540 100.405 286.225 100.545 ;
        RECT 284.540 100.360 284.830 100.405 ;
        RECT 285.905 100.345 286.225 100.405 ;
        RECT 289.140 100.360 289.430 100.590 ;
        RECT 291.440 100.545 291.730 100.590 ;
        RECT 293.725 100.545 294.045 100.605 ;
        RECT 298.325 100.545 298.645 100.605 ;
        RECT 291.440 100.405 294.045 100.545 ;
        RECT 291.440 100.360 291.730 100.405 ;
        RECT 275.320 100.205 275.970 100.250 ;
        RECT 278.920 100.205 279.210 100.250 ;
        RECT 280.385 100.205 280.705 100.265 ;
        RECT 275.320 100.065 280.705 100.205 ;
        RECT 275.320 100.020 275.970 100.065 ;
        RECT 278.620 100.020 279.210 100.065 ;
        RECT 256.555 99.725 258.995 99.865 ;
        RECT 259.700 99.865 259.990 99.910 ;
        RECT 262.445 99.865 262.765 99.925 ;
        RECT 259.700 99.725 262.765 99.865 ;
        RECT 211.845 99.525 212.165 99.585 ;
        RECT 217.840 99.525 218.130 99.570 ;
        RECT 226.105 99.525 226.425 99.585 ;
        RECT 203.655 99.385 211.615 99.525 ;
        RECT 189.270 99.185 189.560 99.230 ;
        RECT 191.160 99.185 191.450 99.230 ;
        RECT 194.280 99.185 194.570 99.230 ;
        RECT 184.795 99.045 185.395 99.185 ;
        RECT 185.255 98.845 185.395 99.045 ;
        RECT 189.270 99.045 194.570 99.185 ;
        RECT 189.270 99.000 189.560 99.045 ;
        RECT 191.160 99.000 191.450 99.045 ;
        RECT 194.280 99.000 194.570 99.045 ;
        RECT 197.600 99.000 197.890 99.230 ;
        RECT 205.980 99.185 206.270 99.230 ;
        RECT 209.100 99.185 209.390 99.230 ;
        RECT 210.990 99.185 211.280 99.230 ;
        RECT 198.135 99.045 205.635 99.185 ;
        RECT 192.065 98.845 192.385 98.905 ;
        RECT 185.255 98.705 192.385 98.845 ;
        RECT 192.065 98.645 192.385 98.705 ;
        RECT 192.985 98.845 193.305 98.905 ;
        RECT 198.135 98.845 198.275 99.045 ;
        RECT 192.985 98.705 198.275 98.845 ;
        RECT 203.120 98.845 203.410 98.890 ;
        RECT 204.945 98.845 205.265 98.905 ;
        RECT 203.120 98.705 205.265 98.845 ;
        RECT 205.495 98.845 205.635 99.045 ;
        RECT 205.980 99.045 211.280 99.185 ;
        RECT 211.475 99.185 211.615 99.385 ;
        RECT 211.845 99.385 226.425 99.525 ;
        RECT 211.845 99.325 212.165 99.385 ;
        RECT 217.840 99.340 218.130 99.385 ;
        RECT 226.105 99.325 226.425 99.385 ;
        RECT 229.325 99.325 229.645 99.585 ;
        RECT 256.555 99.525 256.695 99.725 ;
        RECT 259.700 99.680 259.990 99.725 ;
        RECT 262.445 99.665 262.765 99.725 ;
        RECT 263.825 99.865 264.145 99.925 ;
        RECT 264.760 99.865 265.050 99.910 ;
        RECT 263.825 99.725 265.050 99.865 ;
        RECT 263.825 99.665 264.145 99.725 ;
        RECT 264.760 99.680 265.050 99.725 ;
        RECT 272.125 99.865 272.415 99.910 ;
        RECT 273.960 99.865 274.250 99.910 ;
        RECT 277.540 99.865 277.830 99.910 ;
        RECT 272.125 99.725 277.830 99.865 ;
        RECT 272.125 99.680 272.415 99.725 ;
        RECT 273.960 99.680 274.250 99.725 ;
        RECT 277.540 99.680 277.830 99.725 ;
        RECT 278.620 99.705 278.910 100.020 ;
        RECT 280.385 100.005 280.705 100.065 ;
        RECT 281.305 100.205 281.625 100.265 ;
        RECT 289.215 100.205 289.355 100.360 ;
        RECT 293.725 100.345 294.045 100.405 ;
        RECT 294.275 100.405 298.645 100.545 ;
        RECT 294.275 100.205 294.415 100.405 ;
        RECT 298.325 100.345 298.645 100.405 ;
        RECT 300.625 100.545 300.945 100.605 ;
        RECT 308.000 100.545 308.290 100.590 ;
        RECT 300.625 100.405 308.290 100.545 ;
        RECT 300.625 100.345 300.945 100.405 ;
        RECT 308.000 100.360 308.290 100.405 ;
        RECT 281.305 100.065 289.355 100.205 ;
        RECT 290.135 100.065 294.415 100.205 ;
        RECT 298.785 100.205 299.105 100.265 ;
        RECT 299.700 100.205 300.350 100.250 ;
        RECT 303.300 100.205 303.590 100.250 ;
        RECT 298.785 100.065 303.590 100.205 ;
        RECT 281.305 100.005 281.625 100.065 ;
        RECT 280.845 99.865 281.165 99.925 ;
        RECT 282.240 99.865 282.530 99.910 ;
        RECT 285.445 99.865 285.765 99.925 ;
        RECT 280.845 99.725 285.765 99.865 ;
        RECT 280.845 99.665 281.165 99.725 ;
        RECT 282.240 99.680 282.530 99.725 ;
        RECT 285.445 99.665 285.765 99.725 ;
        RECT 286.365 99.665 286.685 99.925 ;
        RECT 287.745 99.865 288.065 99.925 ;
        RECT 290.135 99.910 290.275 100.065 ;
        RECT 298.785 100.005 299.105 100.065 ;
        RECT 299.700 100.020 300.350 100.065 ;
        RECT 303.000 100.020 303.590 100.065 ;
        RECT 303.845 100.205 304.165 100.265 ;
        RECT 303.845 100.065 307.295 100.205 ;
        RECT 288.220 99.865 288.510 99.910 ;
        RECT 287.745 99.725 288.510 99.865 ;
        RECT 287.745 99.665 288.065 99.725 ;
        RECT 288.220 99.680 288.510 99.725 ;
        RECT 290.060 99.680 290.350 99.910 ;
        RECT 293.280 99.680 293.570 99.910 ;
        RECT 294.645 99.865 294.965 99.925 ;
        RECT 296.040 99.865 296.330 99.910 ;
        RECT 294.645 99.725 296.330 99.865 ;
        RECT 246.895 99.385 256.695 99.525 ;
        RECT 256.925 99.525 257.245 99.585 ;
        RECT 257.860 99.525 258.150 99.570 ;
        RECT 261.985 99.525 262.305 99.585 ;
        RECT 256.925 99.385 262.305 99.525 ;
        RECT 246.895 99.245 247.035 99.385 ;
        RECT 256.925 99.325 257.245 99.385 ;
        RECT 257.860 99.340 258.150 99.385 ;
        RECT 261.985 99.325 262.305 99.385 ;
        RECT 264.285 99.525 264.605 99.585 ;
        RECT 269.345 99.525 269.665 99.585 ;
        RECT 264.285 99.385 269.665 99.525 ;
        RECT 264.285 99.325 264.605 99.385 ;
        RECT 269.345 99.325 269.665 99.385 ;
        RECT 269.820 99.340 270.110 99.570 ;
        RECT 270.265 99.525 270.585 99.585 ;
        RECT 271.660 99.525 271.950 99.570 ;
        RECT 270.265 99.385 271.950 99.525 ;
        RECT 214.145 99.185 214.465 99.245 ;
        RECT 211.475 99.045 214.465 99.185 ;
        RECT 205.980 99.000 206.270 99.045 ;
        RECT 209.100 99.000 209.390 99.045 ;
        RECT 210.990 99.000 211.280 99.045 ;
        RECT 214.145 98.985 214.465 99.045 ;
        RECT 218.710 99.185 219.000 99.230 ;
        RECT 220.600 99.185 220.890 99.230 ;
        RECT 223.720 99.185 224.010 99.230 ;
        RECT 218.710 99.045 224.010 99.185 ;
        RECT 218.710 99.000 219.000 99.045 ;
        RECT 220.600 99.000 220.890 99.045 ;
        RECT 223.720 99.000 224.010 99.045 ;
        RECT 224.265 99.185 224.585 99.245 ;
        RECT 228.880 99.185 229.170 99.230 ;
        RECT 224.265 99.045 229.170 99.185 ;
        RECT 224.265 98.985 224.585 99.045 ;
        RECT 228.880 99.000 229.170 99.045 ;
        RECT 240.790 99.185 241.080 99.230 ;
        RECT 242.680 99.185 242.970 99.230 ;
        RECT 245.800 99.185 246.090 99.230 ;
        RECT 240.790 99.045 246.090 99.185 ;
        RECT 240.790 99.000 241.080 99.045 ;
        RECT 242.680 99.000 242.970 99.045 ;
        RECT 245.800 99.000 246.090 99.045 ;
        RECT 246.805 98.985 247.125 99.245 ;
        RECT 249.990 99.185 250.280 99.230 ;
        RECT 251.880 99.185 252.170 99.230 ;
        RECT 255.000 99.185 255.290 99.230 ;
        RECT 249.990 99.045 255.290 99.185 ;
        RECT 249.990 99.000 250.280 99.045 ;
        RECT 251.880 99.000 252.170 99.045 ;
        RECT 255.000 99.000 255.290 99.045 ;
        RECT 256.465 99.185 256.785 99.245 ;
        RECT 263.840 99.185 264.130 99.230 ;
        RECT 256.465 99.045 264.130 99.185 ;
        RECT 256.465 98.985 256.785 99.045 ;
        RECT 263.840 99.000 264.130 99.045 ;
        RECT 227.945 98.845 228.265 98.905 ;
        RECT 205.495 98.705 228.265 98.845 ;
        RECT 192.985 98.645 193.305 98.705 ;
        RECT 203.120 98.660 203.410 98.705 ;
        RECT 204.945 98.645 205.265 98.705 ;
        RECT 227.945 98.645 228.265 98.705 ;
        RECT 247.725 98.845 248.045 98.905 ;
        RECT 248.660 98.845 248.950 98.890 ;
        RECT 247.725 98.705 248.950 98.845 ;
        RECT 247.725 98.645 248.045 98.705 ;
        RECT 248.660 98.660 248.950 98.705 ;
        RECT 249.105 98.845 249.425 98.905 ;
        RECT 258.305 98.845 258.625 98.905 ;
        RECT 249.105 98.705 258.625 98.845 ;
        RECT 269.895 98.845 270.035 99.340 ;
        RECT 270.265 99.325 270.585 99.385 ;
        RECT 271.660 99.340 271.950 99.385 ;
        RECT 273.025 99.325 273.345 99.585 ;
        RECT 281.320 99.525 281.610 99.570 ;
        RECT 278.175 99.385 281.610 99.525 ;
        RECT 272.530 99.185 272.820 99.230 ;
        RECT 274.420 99.185 274.710 99.230 ;
        RECT 277.540 99.185 277.830 99.230 ;
        RECT 272.530 99.045 277.830 99.185 ;
        RECT 272.530 99.000 272.820 99.045 ;
        RECT 274.420 99.000 274.710 99.045 ;
        RECT 277.540 99.000 277.830 99.045 ;
        RECT 276.705 98.845 277.025 98.905 ;
        RECT 278.175 98.845 278.315 99.385 ;
        RECT 281.320 99.340 281.610 99.385 ;
        RECT 285.905 99.525 286.225 99.585 ;
        RECT 290.135 99.525 290.275 99.680 ;
        RECT 285.905 99.385 290.275 99.525 ;
        RECT 285.905 99.325 286.225 99.385 ;
        RECT 278.545 99.185 278.865 99.245 ;
        RECT 287.300 99.185 287.590 99.230 ;
        RECT 278.545 99.045 287.590 99.185 ;
        RECT 278.545 98.985 278.865 99.045 ;
        RECT 287.300 99.000 287.590 99.045 ;
        RECT 287.745 99.185 288.065 99.245 ;
        RECT 293.355 99.185 293.495 99.680 ;
        RECT 294.645 99.665 294.965 99.725 ;
        RECT 296.040 99.680 296.330 99.725 ;
        RECT 296.505 99.865 296.795 99.910 ;
        RECT 298.340 99.865 298.630 99.910 ;
        RECT 301.920 99.865 302.210 99.910 ;
        RECT 296.505 99.725 302.210 99.865 ;
        RECT 296.505 99.680 296.795 99.725 ;
        RECT 298.340 99.680 298.630 99.725 ;
        RECT 301.920 99.680 302.210 99.725 ;
        RECT 303.000 99.705 303.290 100.020 ;
        RECT 303.845 100.005 304.165 100.065 ;
        RECT 307.155 99.910 307.295 100.065 ;
        RECT 305.240 99.865 305.530 99.910 ;
        RECT 304.165 99.725 305.530 99.865 ;
        RECT 293.725 99.325 294.045 99.585 ;
        RECT 294.185 99.325 294.505 99.585 ;
        RECT 297.420 99.525 297.710 99.570 ;
        RECT 301.085 99.525 301.405 99.585 ;
        RECT 304.165 99.525 304.305 99.725 ;
        RECT 305.240 99.680 305.530 99.725 ;
        RECT 307.080 99.680 307.370 99.910 ;
        RECT 297.420 99.385 301.405 99.525 ;
        RECT 297.420 99.340 297.710 99.385 ;
        RECT 301.085 99.325 301.405 99.385 ;
        RECT 303.015 99.385 304.305 99.525 ;
        RECT 303.015 99.245 303.155 99.385 ;
        RECT 287.745 99.045 293.495 99.185 ;
        RECT 296.910 99.185 297.200 99.230 ;
        RECT 298.800 99.185 299.090 99.230 ;
        RECT 301.920 99.185 302.210 99.230 ;
        RECT 296.910 99.045 302.210 99.185 ;
        RECT 287.745 98.985 288.065 99.045 ;
        RECT 296.910 99.000 297.200 99.045 ;
        RECT 298.800 99.000 299.090 99.045 ;
        RECT 301.920 99.000 302.210 99.045 ;
        RECT 302.925 98.985 303.245 99.245 ;
        RECT 306.160 99.185 306.450 99.230 ;
        RECT 304.395 99.045 306.450 99.185 ;
        RECT 269.895 98.705 278.315 98.845 ;
        RECT 279.005 98.845 279.325 98.905 ;
        RECT 280.400 98.845 280.690 98.890 ;
        RECT 279.005 98.705 280.690 98.845 ;
        RECT 249.105 98.645 249.425 98.705 ;
        RECT 258.305 98.645 258.625 98.705 ;
        RECT 276.705 98.645 277.025 98.705 ;
        RECT 279.005 98.645 279.325 98.705 ;
        RECT 280.400 98.660 280.690 98.705 ;
        RECT 282.685 98.845 283.005 98.905 ;
        RECT 285.460 98.845 285.750 98.890 ;
        RECT 282.685 98.705 285.750 98.845 ;
        RECT 282.685 98.645 283.005 98.705 ;
        RECT 285.460 98.660 285.750 98.705 ;
        RECT 292.805 98.845 293.125 98.905 ;
        RECT 304.395 98.845 304.535 99.045 ;
        RECT 306.160 99.000 306.450 99.045 ;
        RECT 292.805 98.705 304.535 98.845 ;
        RECT 304.780 98.845 305.070 98.890 ;
        RECT 305.685 98.845 306.005 98.905 ;
        RECT 304.780 98.705 306.005 98.845 ;
        RECT 292.805 98.645 293.125 98.705 ;
        RECT 304.780 98.660 305.070 98.705 ;
        RECT 305.685 98.645 306.005 98.705 ;
        RECT 162.095 98.025 311.135 98.505 ;
        RECT 164.480 97.825 164.770 97.870 ;
        RECT 168.145 97.825 168.465 97.885 ;
        RECT 164.480 97.685 168.465 97.825 ;
        RECT 164.480 97.640 164.770 97.685 ;
        RECT 168.145 97.625 168.465 97.685 ;
        RECT 168.605 97.825 168.925 97.885 ;
        RECT 170.920 97.825 171.210 97.870 ;
        RECT 168.605 97.685 171.210 97.825 ;
        RECT 168.605 97.625 168.925 97.685 ;
        RECT 170.920 97.640 171.210 97.685 ;
        RECT 188.845 97.825 189.165 97.885 ;
        RECT 192.080 97.825 192.370 97.870 ;
        RECT 188.845 97.685 192.370 97.825 ;
        RECT 188.845 97.625 189.165 97.685 ;
        RECT 192.080 97.640 192.370 97.685 ;
        RECT 199.900 97.825 200.190 97.870 ;
        RECT 203.105 97.825 203.425 97.885 ;
        RECT 199.900 97.685 203.425 97.825 ;
        RECT 199.900 97.640 200.190 97.685 ;
        RECT 203.105 97.625 203.425 97.685 ;
        RECT 204.025 97.825 204.345 97.885 ;
        RECT 210.465 97.825 210.785 97.885 ;
        RECT 204.025 97.685 210.785 97.825 ;
        RECT 204.025 97.625 204.345 97.685 ;
        RECT 210.465 97.625 210.785 97.685 ;
        RECT 212.320 97.825 212.610 97.870 ;
        RECT 213.685 97.825 214.005 97.885 ;
        RECT 212.320 97.685 214.005 97.825 ;
        RECT 212.320 97.640 212.610 97.685 ;
        RECT 213.685 97.625 214.005 97.685 ;
        RECT 214.145 97.825 214.465 97.885 ;
        RECT 225.185 97.825 225.505 97.885 ;
        RECT 240.840 97.825 241.130 97.870 ;
        RECT 214.145 97.685 225.505 97.825 ;
        RECT 214.145 97.625 214.465 97.685 ;
        RECT 225.185 97.625 225.505 97.685 ;
        RECT 225.735 97.685 241.130 97.825 ;
        RECT 166.320 97.485 166.610 97.530 ;
        RECT 170.445 97.485 170.765 97.545 ;
        RECT 194.365 97.485 194.685 97.545 ;
        RECT 225.735 97.485 225.875 97.685 ;
        RECT 240.840 97.640 241.130 97.685 ;
        RECT 247.265 97.825 247.585 97.885 ;
        RECT 256.925 97.825 257.245 97.885 ;
        RECT 264.285 97.825 264.605 97.885 ;
        RECT 247.265 97.685 257.245 97.825 ;
        RECT 247.265 97.625 247.585 97.685 ;
        RECT 166.320 97.345 170.765 97.485 ;
        RECT 166.320 97.300 166.610 97.345 ;
        RECT 170.445 97.285 170.765 97.345 ;
        RECT 188.015 97.345 194.685 97.485 ;
        RECT 174.140 97.145 174.430 97.190 ;
        RECT 178.740 97.145 179.030 97.190 ;
        RECT 179.645 97.145 179.965 97.205 ;
        RECT 182.880 97.145 183.170 97.190 ;
        RECT 174.140 97.005 183.170 97.145 ;
        RECT 174.140 96.960 174.430 97.005 ;
        RECT 178.740 96.960 179.030 97.005 ;
        RECT 179.645 96.945 179.965 97.005 ;
        RECT 182.880 96.960 183.170 97.005 ;
        RECT 184.720 97.145 185.010 97.190 ;
        RECT 187.465 97.145 187.785 97.205 ;
        RECT 184.720 97.005 187.785 97.145 ;
        RECT 184.720 96.960 185.010 97.005 ;
        RECT 187.465 96.945 187.785 97.005 ;
        RECT 165.385 96.605 165.705 96.865 ;
        RECT 167.240 96.805 167.530 96.850 ;
        RECT 176.425 96.805 176.745 96.865 ;
        RECT 167.240 96.665 176.745 96.805 ;
        RECT 167.240 96.620 167.530 96.665 ;
        RECT 176.425 96.605 176.745 96.665 ;
        RECT 183.800 96.805 184.090 96.850 ;
        RECT 184.245 96.805 184.565 96.865 ;
        RECT 183.800 96.665 184.565 96.805 ;
        RECT 183.800 96.620 184.090 96.665 ;
        RECT 184.245 96.605 184.565 96.665 ;
        RECT 185.180 96.805 185.470 96.850 ;
        RECT 187.005 96.805 187.325 96.865 ;
        RECT 188.015 96.805 188.155 97.345 ;
        RECT 194.365 97.285 194.685 97.345 ;
        RECT 204.115 97.345 225.875 97.485 ;
        RECT 191.160 97.145 191.450 97.190 ;
        RECT 192.065 97.145 192.385 97.205 ;
        RECT 195.300 97.145 195.590 97.190 ;
        RECT 200.345 97.145 200.665 97.205 ;
        RECT 191.160 97.005 200.665 97.145 ;
        RECT 191.160 96.960 191.450 97.005 ;
        RECT 192.065 96.945 192.385 97.005 ;
        RECT 195.300 96.960 195.590 97.005 ;
        RECT 200.345 96.945 200.665 97.005 ;
        RECT 185.180 96.665 188.155 96.805 ;
        RECT 189.780 96.805 190.070 96.850 ;
        RECT 191.605 96.805 191.925 96.865 ;
        RECT 189.780 96.665 191.925 96.805 ;
        RECT 185.180 96.620 185.470 96.665 ;
        RECT 187.005 96.605 187.325 96.665 ;
        RECT 189.780 96.620 190.070 96.665 ;
        RECT 191.605 96.605 191.925 96.665 ;
        RECT 193.920 96.805 194.210 96.850 ;
        RECT 196.205 96.805 196.525 96.865 ;
        RECT 198.965 96.805 199.285 96.865 ;
        RECT 204.115 96.850 204.255 97.345 ;
        RECT 226.120 97.300 226.410 97.530 ;
        RECT 226.565 97.485 226.885 97.545 ;
        RECT 242.665 97.485 242.985 97.545 ;
        RECT 244.505 97.485 244.825 97.545 ;
        RECT 248.200 97.485 248.490 97.530 ;
        RECT 226.565 97.345 244.275 97.485 ;
        RECT 204.945 97.145 205.265 97.205 ;
        RECT 210.005 97.145 210.325 97.205 ;
        RECT 204.945 97.005 209.775 97.145 ;
        RECT 204.945 96.945 205.265 97.005 ;
        RECT 193.920 96.665 199.285 96.805 ;
        RECT 193.920 96.620 194.210 96.665 ;
        RECT 196.205 96.605 196.525 96.665 ;
        RECT 198.965 96.605 199.285 96.665 ;
        RECT 204.040 96.620 204.330 96.850 ;
        RECT 205.420 96.805 205.710 96.850 ;
        RECT 206.325 96.805 206.645 96.865 ;
        RECT 205.420 96.665 206.645 96.805 ;
        RECT 205.420 96.620 205.710 96.665 ;
        RECT 206.325 96.605 206.645 96.665 ;
        RECT 206.785 96.605 207.105 96.865 ;
        RECT 207.705 96.605 208.025 96.865 ;
        RECT 208.625 96.605 208.945 96.865 ;
        RECT 209.635 96.850 209.775 97.005 ;
        RECT 210.005 97.005 225.875 97.145 ;
        RECT 210.005 96.945 210.325 97.005 ;
        RECT 209.560 96.805 209.850 96.850 ;
        RECT 217.825 96.805 218.145 96.865 ;
        RECT 223.360 96.805 223.650 96.850 ;
        RECT 209.560 96.665 223.650 96.805 ;
        RECT 209.560 96.620 209.850 96.665 ;
        RECT 217.825 96.605 218.145 96.665 ;
        RECT 223.360 96.620 223.650 96.665 ;
        RECT 225.185 96.605 225.505 96.865 ;
        RECT 172.760 96.465 173.050 96.510 ;
        RECT 176.885 96.465 177.205 96.525 ;
        RECT 172.760 96.325 177.205 96.465 ;
        RECT 172.760 96.280 173.050 96.325 ;
        RECT 176.885 96.265 177.205 96.325 ;
        RECT 177.360 96.465 177.650 96.510 ;
        RECT 180.105 96.465 180.425 96.525 ;
        RECT 177.360 96.325 180.425 96.465 ;
        RECT 177.360 96.280 177.650 96.325 ;
        RECT 180.105 96.265 180.425 96.325 ;
        RECT 185.625 96.465 185.945 96.525 ;
        RECT 207.260 96.465 207.550 96.510 ;
        RECT 185.625 96.325 207.550 96.465 ;
        RECT 185.625 96.265 185.945 96.325 ;
        RECT 207.260 96.280 207.550 96.325 ;
        RECT 223.805 96.465 224.125 96.525 ;
        RECT 224.280 96.465 224.570 96.510 ;
        RECT 223.805 96.325 224.570 96.465 ;
        RECT 173.220 96.125 173.510 96.170 ;
        RECT 175.045 96.125 175.365 96.185 ;
        RECT 173.220 95.985 175.365 96.125 ;
        RECT 173.220 95.940 173.510 95.985 ;
        RECT 175.045 95.925 175.365 95.985 ;
        RECT 175.505 95.925 175.825 96.185 ;
        RECT 177.820 96.125 178.110 96.170 ;
        RECT 179.645 96.125 179.965 96.185 ;
        RECT 186.085 96.125 186.405 96.185 ;
        RECT 177.820 95.985 186.405 96.125 ;
        RECT 177.820 95.940 178.110 95.985 ;
        RECT 179.645 95.925 179.965 95.985 ;
        RECT 186.085 95.925 186.405 95.985 ;
        RECT 187.925 95.925 188.245 96.185 ;
        RECT 190.225 95.925 190.545 96.185 ;
        RECT 194.380 96.125 194.670 96.170 ;
        RECT 194.825 96.125 195.145 96.185 ;
        RECT 194.380 95.985 195.145 96.125 ;
        RECT 194.380 95.940 194.670 95.985 ;
        RECT 194.825 95.925 195.145 95.985 ;
        RECT 200.345 96.125 200.665 96.185 ;
        RECT 203.120 96.125 203.410 96.170 ;
        RECT 200.345 95.985 203.410 96.125 ;
        RECT 200.345 95.925 200.665 95.985 ;
        RECT 203.120 95.940 203.410 95.985 ;
        RECT 204.945 95.925 205.265 96.185 ;
        RECT 205.880 96.125 206.170 96.170 ;
        RECT 206.785 96.125 207.105 96.185 ;
        RECT 205.880 95.985 207.105 96.125 ;
        RECT 207.335 96.125 207.475 96.280 ;
        RECT 223.805 96.265 224.125 96.325 ;
        RECT 224.280 96.280 224.570 96.325 ;
        RECT 224.740 96.280 225.030 96.510 ;
        RECT 225.735 96.465 225.875 97.005 ;
        RECT 226.195 96.805 226.335 97.300 ;
        RECT 226.565 97.285 226.885 97.345 ;
        RECT 242.665 97.285 242.985 97.345 ;
        RECT 229.415 97.005 243.815 97.145 ;
        RECT 227.500 96.805 227.790 96.850 ;
        RECT 226.195 96.665 227.790 96.805 ;
        RECT 227.500 96.620 227.790 96.665 ;
        RECT 227.945 96.805 228.265 96.865 ;
        RECT 229.415 96.850 229.555 97.005 ;
        RECT 243.675 96.865 243.815 97.005 ;
        RECT 227.945 96.665 228.460 96.805 ;
        RECT 227.945 96.605 228.265 96.665 ;
        RECT 229.340 96.620 229.630 96.850 ;
        RECT 230.030 96.805 230.320 96.850 ;
        RECT 231.625 96.805 231.945 96.865 ;
        RECT 230.030 96.665 231.945 96.805 ;
        RECT 230.030 96.620 230.320 96.665 ;
        RECT 231.625 96.605 231.945 96.665 ;
        RECT 241.745 96.605 242.065 96.865 ;
        RECT 242.220 96.805 242.510 96.850 ;
        RECT 242.220 96.665 243.355 96.805 ;
        RECT 242.220 96.620 242.510 96.665 ;
        RECT 228.880 96.465 229.170 96.510 ;
        RECT 232.085 96.465 232.405 96.525 ;
        RECT 225.735 96.325 232.405 96.465 ;
        RECT 228.880 96.280 229.170 96.325 ;
        RECT 208.625 96.125 208.945 96.185 ;
        RECT 207.335 95.985 208.945 96.125 ;
        RECT 224.815 96.125 224.955 96.280 ;
        RECT 232.085 96.265 232.405 96.325 ;
        RECT 233.925 96.465 234.245 96.525 ;
        RECT 241.285 96.465 241.605 96.525 ;
        RECT 242.680 96.465 242.970 96.510 ;
        RECT 233.925 96.325 242.970 96.465 ;
        RECT 243.215 96.465 243.355 96.665 ;
        RECT 243.585 96.605 243.905 96.865 ;
        RECT 244.135 96.850 244.275 97.345 ;
        RECT 244.505 97.345 248.490 97.485 ;
        RECT 244.505 97.285 244.825 97.345 ;
        RECT 248.200 97.300 248.490 97.345 ;
        RECT 249.105 97.285 249.425 97.545 ;
        RECT 244.060 96.620 244.350 96.850 ;
        RECT 245.900 96.805 246.190 96.850 ;
        RECT 246.805 96.805 247.125 96.865 ;
        RECT 249.170 96.850 249.310 97.285 ;
        RECT 249.655 96.850 249.795 97.685 ;
        RECT 256.925 97.625 257.245 97.685 ;
        RECT 257.475 97.685 264.605 97.825 ;
        RECT 252.800 97.300 253.090 97.530 ;
        RECT 254.625 97.485 254.945 97.545 ;
        RECT 257.475 97.485 257.615 97.685 ;
        RECT 264.285 97.625 264.605 97.685 ;
        RECT 265.205 97.825 265.525 97.885 ;
        RECT 271.660 97.825 271.950 97.870 ;
        RECT 265.205 97.685 271.950 97.825 ;
        RECT 265.205 97.625 265.525 97.685 ;
        RECT 271.660 97.640 271.950 97.685 ;
        RECT 273.025 97.825 273.345 97.885 ;
        RECT 273.960 97.825 274.250 97.870 ;
        RECT 273.025 97.685 274.250 97.825 ;
        RECT 273.025 97.625 273.345 97.685 ;
        RECT 273.960 97.640 274.250 97.685 ;
        RECT 282.225 97.625 282.545 97.885 ;
        RECT 283.605 97.825 283.925 97.885 ;
        RECT 286.380 97.825 286.670 97.870 ;
        RECT 283.605 97.685 286.670 97.825 ;
        RECT 283.605 97.625 283.925 97.685 ;
        RECT 286.380 97.640 286.670 97.685 ;
        RECT 288.205 97.825 288.525 97.885 ;
        RECT 289.600 97.825 289.890 97.870 ;
        RECT 288.205 97.685 289.890 97.825 ;
        RECT 288.205 97.625 288.525 97.685 ;
        RECT 289.600 97.640 289.890 97.685 ;
        RECT 294.185 97.825 294.505 97.885 ;
        RECT 297.865 97.825 298.185 97.885 ;
        RECT 294.185 97.685 298.185 97.825 ;
        RECT 294.185 97.625 294.505 97.685 ;
        RECT 297.865 97.625 298.185 97.685 ;
        RECT 298.325 97.825 298.645 97.885 ;
        RECT 303.400 97.825 303.690 97.870 ;
        RECT 298.325 97.685 303.690 97.825 ;
        RECT 298.325 97.625 298.645 97.685 ;
        RECT 303.400 97.640 303.690 97.685 ;
        RECT 254.625 97.345 257.615 97.485 ;
        RECT 257.860 97.485 258.150 97.530 ;
        RECT 260.145 97.485 260.465 97.545 ;
        RECT 257.860 97.345 260.465 97.485 ;
        RECT 244.595 96.665 245.655 96.805 ;
        RECT 244.595 96.465 244.735 96.665 ;
        RECT 245.515 96.510 245.655 96.665 ;
        RECT 245.900 96.665 247.125 96.805 ;
        RECT 245.900 96.620 246.190 96.665 ;
        RECT 246.805 96.605 247.125 96.665 ;
        RECT 249.095 96.620 249.385 96.850 ;
        RECT 249.580 96.620 249.870 96.850 ;
        RECT 250.025 96.605 250.345 96.865 ;
        RECT 250.955 96.620 251.245 96.850 ;
        RECT 251.420 96.805 251.710 96.850 ;
        RECT 252.875 96.805 253.015 97.300 ;
        RECT 254.625 97.285 254.945 97.345 ;
        RECT 257.860 97.300 258.150 97.345 ;
        RECT 260.145 97.285 260.465 97.345 ;
        RECT 262.905 97.485 263.225 97.545 ;
        RECT 269.820 97.485 270.110 97.530 ;
        RECT 285.905 97.485 286.225 97.545 ;
        RECT 262.905 97.345 270.110 97.485 ;
        RECT 262.905 97.285 263.225 97.345 ;
        RECT 269.820 97.300 270.110 97.345 ;
        RECT 275.875 97.345 286.225 97.485 ;
        RECT 275.325 97.145 275.645 97.205 ;
        RECT 251.420 96.665 253.015 96.805 ;
        RECT 253.335 97.005 275.645 97.145 ;
        RECT 251.420 96.620 251.710 96.665 ;
        RECT 243.215 96.325 244.735 96.465 ;
        RECT 233.925 96.265 234.245 96.325 ;
        RECT 241.285 96.265 241.605 96.325 ;
        RECT 242.680 96.280 242.970 96.325 ;
        RECT 244.980 96.280 245.270 96.510 ;
        RECT 245.440 96.465 245.730 96.510 ;
        RECT 248.185 96.465 248.505 96.525 ;
        RECT 245.440 96.325 248.505 96.465 ;
        RECT 251.030 96.465 251.170 96.620 ;
        RECT 251.865 96.465 252.185 96.525 ;
        RECT 253.335 96.465 253.475 97.005 ;
        RECT 253.705 96.605 254.025 96.865 ;
        RECT 254.165 96.605 254.485 96.865 ;
        RECT 255.560 96.620 255.850 96.850 ;
        RECT 256.020 96.805 256.310 96.850 ;
        RECT 257.385 96.805 257.705 96.865 ;
        RECT 256.020 96.665 257.705 96.805 ;
        RECT 256.020 96.620 256.310 96.665 ;
        RECT 251.030 96.325 253.475 96.465 ;
        RECT 245.440 96.280 245.730 96.325 ;
        RECT 227.485 96.125 227.805 96.185 ;
        RECT 224.815 95.985 227.805 96.125 ;
        RECT 205.880 95.940 206.170 95.985 ;
        RECT 206.785 95.925 207.105 95.985 ;
        RECT 208.625 95.925 208.945 95.985 ;
        RECT 227.485 95.925 227.805 95.985 ;
        RECT 228.405 96.125 228.725 96.185 ;
        RECT 230.720 96.125 231.010 96.170 ;
        RECT 228.405 95.985 231.010 96.125 ;
        RECT 228.405 95.925 228.725 95.985 ;
        RECT 230.720 95.940 231.010 95.985 ;
        RECT 232.545 96.125 232.865 96.185 ;
        RECT 245.055 96.125 245.195 96.280 ;
        RECT 248.185 96.265 248.505 96.325 ;
        RECT 251.865 96.265 252.185 96.325 ;
        RECT 254.625 96.265 254.945 96.525 ;
        RECT 255.635 96.465 255.775 96.620 ;
        RECT 257.385 96.605 257.705 96.665 ;
        RECT 257.860 96.805 258.150 96.850 ;
        RECT 258.305 96.805 258.625 96.865 ;
        RECT 257.860 96.665 258.625 96.805 ;
        RECT 257.860 96.620 258.150 96.665 ;
        RECT 258.305 96.605 258.625 96.665 ;
        RECT 258.765 96.605 259.085 96.865 ;
        RECT 270.815 96.850 270.955 97.005 ;
        RECT 275.325 96.945 275.645 97.005 ;
        RECT 270.740 96.620 271.030 96.850 ;
        RECT 272.565 96.605 272.885 96.865 ;
        RECT 275.875 96.805 276.015 97.345 ;
        RECT 285.905 97.285 286.225 97.345 ;
        RECT 286.825 97.485 287.145 97.545 ;
        RECT 290.980 97.485 291.270 97.530 ;
        RECT 286.825 97.345 291.270 97.485 ;
        RECT 286.825 97.285 287.145 97.345 ;
        RECT 290.980 97.300 291.270 97.345 ;
        RECT 295.530 97.485 295.820 97.530 ;
        RECT 297.420 97.485 297.710 97.530 ;
        RECT 300.540 97.485 300.830 97.530 ;
        RECT 295.530 97.345 300.830 97.485 ;
        RECT 295.530 97.300 295.820 97.345 ;
        RECT 297.420 97.300 297.710 97.345 ;
        RECT 300.540 97.300 300.830 97.345 ;
        RECT 301.085 97.485 301.405 97.545 ;
        RECT 304.320 97.485 304.610 97.530 ;
        RECT 301.085 97.345 304.610 97.485 ;
        RECT 301.085 97.285 301.405 97.345 ;
        RECT 304.320 97.300 304.610 97.345 ;
        RECT 276.705 97.145 277.025 97.205 ;
        RECT 279.020 97.145 279.310 97.190 ;
        RECT 279.465 97.145 279.785 97.205 ;
        RECT 276.705 97.005 279.785 97.145 ;
        RECT 276.705 96.945 277.025 97.005 ;
        RECT 279.020 96.960 279.310 97.005 ;
        RECT 279.465 96.945 279.785 97.005 ;
        RECT 279.925 96.945 280.245 97.205 ;
        RECT 283.160 97.145 283.450 97.190 ;
        RECT 283.605 97.145 283.925 97.205 ;
        RECT 283.160 97.005 283.925 97.145 ;
        RECT 283.160 96.960 283.450 97.005 ;
        RECT 283.605 96.945 283.925 97.005 ;
        RECT 285.000 97.145 285.290 97.190 ;
        RECT 294.185 97.145 294.505 97.205 ;
        RECT 285.000 97.005 294.505 97.145 ;
        RECT 285.000 96.960 285.290 97.005 ;
        RECT 294.185 96.945 294.505 97.005 ;
        RECT 294.645 97.145 294.965 97.205 ;
        RECT 296.025 97.145 296.345 97.205 ;
        RECT 294.645 97.005 296.345 97.145 ;
        RECT 294.645 96.945 294.965 97.005 ;
        RECT 296.025 96.945 296.345 97.005 ;
        RECT 299.705 97.145 300.025 97.205 ;
        RECT 307.080 97.145 307.370 97.190 ;
        RECT 299.705 97.005 307.370 97.145 ;
        RECT 299.705 96.945 300.025 97.005 ;
        RECT 307.080 96.960 307.370 97.005 ;
        RECT 274.955 96.665 276.015 96.805 ;
        RECT 274.955 96.465 275.095 96.665 ;
        RECT 276.245 96.605 276.565 96.865 ;
        RECT 277.165 96.805 277.485 96.865 ;
        RECT 280.400 96.805 280.690 96.850 ;
        RECT 277.165 96.665 280.690 96.805 ;
        RECT 277.165 96.605 277.485 96.665 ;
        RECT 280.400 96.620 280.690 96.665 ;
        RECT 282.685 96.605 283.005 96.865 ;
        RECT 284.080 96.620 284.370 96.850 ;
        RECT 284.525 96.805 284.845 96.865 ;
        RECT 285.460 96.805 285.750 96.850 ;
        RECT 284.525 96.665 285.750 96.805 ;
        RECT 278.545 96.465 278.865 96.525 ;
        RECT 283.145 96.465 283.465 96.525 ;
        RECT 284.155 96.465 284.295 96.620 ;
        RECT 284.525 96.605 284.845 96.665 ;
        RECT 285.460 96.620 285.750 96.665 ;
        RECT 288.665 96.605 288.985 96.865 ;
        RECT 291.900 96.805 292.190 96.850 ;
        RECT 292.805 96.805 293.125 96.865 ;
        RECT 291.900 96.665 293.125 96.805 ;
        RECT 291.900 96.620 292.190 96.665 ;
        RECT 292.805 96.605 293.125 96.665 ;
        RECT 295.125 96.805 295.415 96.850 ;
        RECT 296.960 96.805 297.250 96.850 ;
        RECT 300.540 96.805 300.830 96.850 ;
        RECT 295.125 96.665 300.830 96.805 ;
        RECT 295.125 96.620 295.415 96.665 ;
        RECT 296.960 96.620 297.250 96.665 ;
        RECT 300.540 96.620 300.830 96.665 ;
        RECT 301.620 96.805 301.910 96.825 ;
        RECT 305.225 96.805 305.545 96.865 ;
        RECT 301.620 96.665 305.545 96.805 ;
        RECT 255.635 96.325 275.095 96.465 ;
        RECT 275.415 96.325 284.295 96.465 ;
        RECT 296.040 96.465 296.330 96.510 ;
        RECT 296.485 96.465 296.805 96.525 ;
        RECT 301.620 96.510 301.910 96.665 ;
        RECT 305.225 96.605 305.545 96.665 ;
        RECT 296.040 96.325 296.805 96.465 ;
        RECT 232.545 95.985 245.195 96.125 ;
        RECT 246.345 96.125 246.665 96.185 ;
        RECT 246.820 96.125 247.110 96.170 ;
        RECT 246.345 95.985 247.110 96.125 ;
        RECT 232.545 95.925 232.865 95.985 ;
        RECT 246.345 95.925 246.665 95.985 ;
        RECT 246.820 95.940 247.110 95.985 ;
        RECT 248.645 96.125 248.965 96.185 ;
        RECT 255.865 96.125 256.005 96.325 ;
        RECT 248.645 95.985 256.005 96.125 ;
        RECT 257.845 96.125 258.165 96.185 ;
        RECT 275.415 96.125 275.555 96.325 ;
        RECT 278.545 96.265 278.865 96.325 ;
        RECT 283.145 96.265 283.465 96.325 ;
        RECT 296.040 96.280 296.330 96.325 ;
        RECT 296.485 96.265 296.805 96.325 ;
        RECT 298.320 96.465 298.970 96.510 ;
        RECT 301.620 96.465 302.210 96.510 ;
        RECT 306.620 96.465 306.910 96.510 ;
        RECT 307.065 96.465 307.385 96.525 ;
        RECT 298.320 96.325 302.210 96.465 ;
        RECT 298.320 96.280 298.970 96.325 ;
        RECT 301.920 96.280 302.210 96.325 ;
        RECT 302.555 96.325 307.385 96.465 ;
        RECT 257.845 95.985 275.555 96.125 ;
        RECT 275.785 96.125 276.105 96.185 ;
        RECT 279.005 96.125 279.325 96.185 ;
        RECT 275.785 95.985 279.325 96.125 ;
        RECT 248.645 95.925 248.965 95.985 ;
        RECT 257.845 95.925 258.165 95.985 ;
        RECT 275.785 95.925 276.105 95.985 ;
        RECT 279.005 95.925 279.325 95.985 ;
        RECT 279.925 96.125 280.245 96.185 ;
        RECT 302.555 96.125 302.695 96.325 ;
        RECT 306.620 96.280 306.910 96.325 ;
        RECT 307.065 96.265 307.385 96.325 ;
        RECT 279.925 95.985 302.695 96.125 ;
        RECT 279.925 95.925 280.245 95.985 ;
        RECT 306.145 95.925 306.465 96.185 ;
        RECT 162.095 95.305 311.135 95.785 ;
        RECT 179.200 95.105 179.490 95.150 ;
        RECT 180.105 95.105 180.425 95.165 ;
        RECT 185.625 95.105 185.945 95.165 ;
        RECT 179.200 94.965 185.945 95.105 ;
        RECT 179.200 94.920 179.490 94.965 ;
        RECT 180.105 94.905 180.425 94.965 ;
        RECT 185.625 94.905 185.945 94.965 ;
        RECT 191.145 94.905 191.465 95.165 ;
        RECT 192.065 94.905 192.385 95.165 ;
        RECT 207.720 95.105 208.010 95.150 ;
        RECT 208.165 95.105 208.485 95.165 ;
        RECT 210.005 95.105 210.325 95.165 ;
        RECT 207.720 94.965 210.325 95.105 ;
        RECT 207.720 94.920 208.010 94.965 ;
        RECT 208.165 94.905 208.485 94.965 ;
        RECT 210.005 94.905 210.325 94.965 ;
        RECT 215.065 95.105 215.385 95.165 ;
        RECT 226.120 95.105 226.410 95.150 ;
        RECT 215.065 94.965 226.410 95.105 ;
        RECT 215.065 94.905 215.385 94.965 ;
        RECT 226.120 94.920 226.410 94.965 ;
        RECT 227.945 94.905 228.265 95.165 ;
        RECT 231.625 95.105 231.945 95.165 ;
        RECT 231.625 94.965 235.995 95.105 ;
        RECT 231.625 94.905 231.945 94.965 ;
        RECT 169.985 94.765 170.305 94.825 ;
        RECT 172.285 94.765 172.605 94.825 ;
        RECT 174.120 94.765 174.770 94.810 ;
        RECT 177.720 94.765 178.010 94.810 ;
        RECT 169.985 94.625 178.010 94.765 ;
        RECT 169.985 94.565 170.305 94.625 ;
        RECT 172.285 94.565 172.605 94.625 ;
        RECT 174.120 94.580 174.770 94.625 ;
        RECT 177.420 94.580 178.010 94.625 ;
        RECT 189.780 94.765 190.070 94.810 ;
        RECT 192.525 94.765 192.845 94.825 ;
        RECT 223.345 94.765 223.665 94.825 ;
        RECT 189.780 94.625 192.845 94.765 ;
        RECT 189.780 94.580 190.070 94.625 ;
        RECT 164.925 94.225 165.245 94.485 ;
        RECT 167.225 94.425 167.545 94.485 ;
        RECT 170.460 94.425 170.750 94.470 ;
        RECT 167.225 94.285 170.750 94.425 ;
        RECT 167.225 94.225 167.545 94.285 ;
        RECT 170.460 94.240 170.750 94.285 ;
        RECT 170.925 94.425 171.215 94.470 ;
        RECT 172.760 94.425 173.050 94.470 ;
        RECT 176.340 94.425 176.630 94.470 ;
        RECT 170.925 94.285 176.630 94.425 ;
        RECT 170.925 94.240 171.215 94.285 ;
        RECT 172.760 94.240 173.050 94.285 ;
        RECT 176.340 94.240 176.630 94.285 ;
        RECT 177.420 94.265 177.710 94.580 ;
        RECT 192.525 94.565 192.845 94.625 ;
        RECT 208.255 94.625 223.665 94.765 ;
        RECT 184.245 94.425 184.565 94.485 ;
        RECT 189.305 94.425 189.625 94.485 ;
        RECT 192.985 94.425 193.305 94.485 ;
        RECT 184.245 94.285 193.305 94.425 ;
        RECT 184.245 94.225 184.565 94.285 ;
        RECT 189.305 94.225 189.625 94.285 ;
        RECT 192.985 94.225 193.305 94.285 ;
        RECT 193.920 94.425 194.210 94.470 ;
        RECT 204.025 94.425 204.345 94.485 ;
        RECT 193.920 94.285 204.345 94.425 ;
        RECT 193.920 94.240 194.210 94.285 ;
        RECT 204.025 94.225 204.345 94.285 ;
        RECT 206.785 94.225 207.105 94.485 ;
        RECT 208.255 94.470 208.395 94.625 ;
        RECT 223.345 94.565 223.665 94.625 ;
        RECT 227.500 94.765 227.790 94.810 ;
        RECT 228.035 94.765 228.175 94.905 ;
        RECT 235.305 94.765 235.625 94.825 ;
        RECT 227.500 94.625 228.175 94.765 ;
        RECT 228.955 94.625 235.625 94.765 ;
        RECT 235.855 94.765 235.995 94.965 ;
        RECT 241.835 94.965 249.795 95.105 ;
        RECT 241.835 94.765 241.975 94.965 ;
        RECT 235.855 94.625 241.975 94.765 ;
        RECT 227.500 94.580 227.790 94.625 ;
        RECT 208.180 94.240 208.470 94.470 ;
        RECT 208.625 94.225 208.945 94.485 ;
        RECT 209.545 94.225 209.865 94.485 ;
        RECT 210.005 94.225 210.325 94.485 ;
        RECT 210.465 94.425 210.785 94.485 ;
        RECT 226.565 94.470 226.885 94.485 ;
        RECT 210.465 94.285 225.415 94.425 ;
        RECT 210.465 94.225 210.785 94.285 ;
        RECT 171.840 94.085 172.130 94.130 ;
        RECT 175.505 94.085 175.825 94.145 ;
        RECT 171.840 93.945 175.825 94.085 ;
        RECT 171.840 93.900 172.130 93.945 ;
        RECT 175.505 93.885 175.825 93.945 ;
        RECT 194.365 93.885 194.685 94.145 ;
        RECT 203.105 94.085 203.425 94.145 ;
        RECT 209.635 94.085 209.775 94.225 ;
        RECT 203.105 93.945 209.775 94.085 ;
        RECT 203.105 93.885 203.425 93.945 ;
        RECT 171.330 93.745 171.620 93.790 ;
        RECT 173.220 93.745 173.510 93.790 ;
        RECT 176.340 93.745 176.630 93.790 ;
        RECT 171.330 93.605 176.630 93.745 ;
        RECT 171.330 93.560 171.620 93.605 ;
        RECT 173.220 93.560 173.510 93.605 ;
        RECT 176.340 93.560 176.630 93.605 ;
        RECT 198.965 93.745 199.285 93.805 ;
        RECT 224.725 93.745 225.045 93.805 ;
        RECT 198.965 93.605 225.045 93.745 ;
        RECT 225.275 93.745 225.415 94.285 ;
        RECT 226.565 94.240 227.100 94.470 ;
        RECT 226.565 94.225 226.885 94.240 ;
        RECT 227.945 94.225 228.265 94.485 ;
        RECT 228.955 94.470 229.095 94.625 ;
        RECT 235.305 94.565 235.625 94.625 ;
        RECT 242.665 94.565 242.985 94.825 ;
        RECT 243.140 94.765 243.430 94.810 ;
        RECT 243.140 94.625 248.415 94.765 ;
        RECT 243.140 94.580 243.430 94.625 ;
        RECT 228.875 94.425 229.165 94.470 ;
        RECT 228.495 94.285 229.165 94.425 ;
        RECT 227.485 94.085 227.805 94.145 ;
        RECT 228.495 94.085 228.635 94.285 ;
        RECT 228.875 94.240 229.165 94.285 ;
        RECT 229.340 94.425 229.630 94.470 ;
        RECT 242.195 94.425 242.485 94.470 ;
        RECT 229.340 94.285 241.515 94.425 ;
        RECT 229.340 94.240 229.630 94.285 ;
        RECT 227.485 93.945 228.635 94.085 ;
        RECT 227.485 93.885 227.805 93.945 ;
        RECT 232.545 93.745 232.865 93.805 ;
        RECT 241.375 93.790 241.515 94.285 ;
        RECT 242.195 94.285 242.895 94.425 ;
        RECT 242.195 94.240 242.485 94.285 ;
        RECT 242.755 94.145 242.895 94.285 ;
        RECT 244.055 94.240 244.345 94.470 ;
        RECT 244.520 94.425 244.810 94.470 ;
        RECT 246.820 94.425 247.110 94.470 ;
        RECT 244.520 94.285 247.110 94.425 ;
        RECT 244.520 94.240 244.810 94.285 ;
        RECT 246.820 94.240 247.110 94.285 ;
        RECT 247.265 94.425 247.585 94.485 ;
        RECT 248.275 94.470 248.415 94.625 ;
        RECT 248.645 94.565 248.965 94.825 ;
        RECT 249.105 94.470 249.425 94.485 ;
        RECT 247.265 94.285 247.780 94.425 ;
        RECT 242.665 93.885 242.985 94.145 ;
        RECT 244.135 94.085 244.275 94.240 ;
        RECT 244.965 94.085 245.285 94.145 ;
        RECT 245.885 94.085 246.205 94.145 ;
        RECT 244.135 93.945 246.205 94.085 ;
        RECT 244.965 93.885 245.285 93.945 ;
        RECT 245.885 93.885 246.205 93.945 ;
        RECT 225.275 93.605 232.865 93.745 ;
        RECT 198.965 93.545 199.285 93.605 ;
        RECT 224.725 93.545 225.045 93.605 ;
        RECT 232.545 93.545 232.865 93.605 ;
        RECT 241.300 93.560 241.590 93.790 ;
        RECT 164.005 93.205 164.325 93.465 ;
        RECT 186.085 93.405 186.405 93.465 ;
        RECT 194.825 93.405 195.145 93.465 ;
        RECT 186.085 93.265 195.145 93.405 ;
        RECT 186.085 93.205 186.405 93.265 ;
        RECT 194.825 93.205 195.145 93.265 ;
        RECT 205.865 93.205 206.185 93.465 ;
        RECT 211.400 93.405 211.690 93.450 ;
        RECT 214.145 93.405 214.465 93.465 ;
        RECT 211.400 93.265 214.465 93.405 ;
        RECT 211.400 93.220 211.690 93.265 ;
        RECT 214.145 93.205 214.465 93.265 ;
        RECT 216.905 93.405 217.225 93.465 ;
        RECT 225.645 93.405 225.965 93.465 ;
        RECT 227.485 93.405 227.805 93.465 ;
        RECT 216.905 93.265 227.805 93.405 ;
        RECT 216.905 93.205 217.225 93.265 ;
        RECT 225.645 93.205 225.965 93.265 ;
        RECT 227.485 93.205 227.805 93.265 ;
        RECT 227.945 93.405 228.265 93.465 ;
        RECT 233.925 93.405 234.245 93.465 ;
        RECT 227.945 93.265 234.245 93.405 ;
        RECT 227.945 93.205 228.265 93.265 ;
        RECT 233.925 93.205 234.245 93.265 ;
        RECT 241.745 93.405 242.065 93.465 ;
        RECT 245.885 93.405 246.205 93.465 ;
        RECT 241.745 93.265 246.205 93.405 ;
        RECT 246.895 93.405 247.035 94.240 ;
        RECT 247.265 94.225 247.585 94.285 ;
        RECT 248.200 94.240 248.490 94.470 ;
        RECT 249.105 94.425 249.435 94.470 ;
        RECT 248.935 94.285 249.435 94.425 ;
        RECT 249.655 94.425 249.795 94.965 ;
        RECT 250.040 94.920 250.330 95.150 ;
        RECT 250.485 95.105 250.805 95.165 ;
        RECT 263.825 95.105 264.145 95.165 ;
        RECT 277.625 95.105 277.945 95.165 ;
        RECT 250.485 94.965 254.395 95.105 ;
        RECT 250.115 94.765 250.255 94.920 ;
        RECT 250.485 94.905 250.805 94.965 ;
        RECT 250.115 94.625 253.935 94.765 ;
        RECT 251.405 94.470 251.725 94.485 ;
        RECT 251.395 94.425 251.725 94.470 ;
        RECT 249.655 94.285 250.715 94.425 ;
        RECT 251.210 94.285 251.725 94.425 ;
        RECT 249.105 94.240 249.435 94.285 ;
        RECT 248.275 94.085 248.415 94.240 ;
        RECT 249.105 94.225 249.425 94.240 ;
        RECT 248.645 94.085 248.965 94.145 ;
        RECT 248.275 93.945 248.965 94.085 ;
        RECT 250.575 94.085 250.715 94.285 ;
        RECT 251.395 94.240 251.725 94.285 ;
        RECT 251.405 94.225 251.725 94.240 ;
        RECT 251.865 94.225 252.185 94.485 ;
        RECT 252.325 94.225 252.645 94.485 ;
        RECT 252.785 94.470 253.105 94.485 ;
        RECT 253.795 94.470 253.935 94.625 ;
        RECT 252.785 94.240 253.270 94.470 ;
        RECT 253.720 94.240 254.010 94.470 ;
        RECT 254.255 94.425 254.395 94.965 ;
        RECT 263.825 94.965 277.945 95.105 ;
        RECT 263.825 94.905 264.145 94.965 ;
        RECT 277.625 94.905 277.945 94.965 ;
        RECT 279.465 94.905 279.785 95.165 ;
        RECT 293.725 94.905 294.045 95.165 ;
        RECT 296.500 95.105 296.790 95.150 ;
        RECT 296.945 95.105 297.265 95.165 ;
        RECT 296.500 94.965 297.265 95.105 ;
        RECT 296.500 94.920 296.790 94.965 ;
        RECT 296.945 94.905 297.265 94.965 ;
        RECT 298.340 95.105 298.630 95.150 ;
        RECT 298.785 95.105 299.105 95.165 ;
        RECT 298.340 94.965 299.105 95.105 ;
        RECT 298.340 94.920 298.630 94.965 ;
        RECT 298.785 94.905 299.105 94.965 ;
        RECT 300.640 94.920 300.930 95.150 ;
        RECT 304.765 95.105 305.085 95.165 ;
        RECT 305.700 95.105 305.990 95.150 ;
        RECT 304.765 94.965 305.990 95.105 ;
        RECT 255.085 94.765 255.405 94.825 ;
        RECT 280.845 94.765 281.165 94.825 ;
        RECT 255.085 94.625 281.165 94.765 ;
        RECT 255.085 94.565 255.405 94.625 ;
        RECT 276.705 94.425 277.025 94.485 ;
        RECT 254.255 94.285 277.025 94.425 ;
        RECT 252.785 94.225 253.105 94.240 ;
        RECT 276.705 94.225 277.025 94.285 ;
        RECT 277.165 94.225 277.485 94.485 ;
        RECT 277.715 94.470 277.855 94.625 ;
        RECT 280.845 94.565 281.165 94.625 ;
        RECT 285.445 94.765 285.765 94.825 ;
        RECT 295.565 94.765 295.885 94.825 ;
        RECT 300.715 94.765 300.855 94.920 ;
        RECT 304.765 94.905 305.085 94.965 ;
        RECT 305.700 94.920 305.990 94.965 ;
        RECT 306.605 95.105 306.925 95.165 ;
        RECT 308.000 95.105 308.290 95.150 ;
        RECT 306.605 94.965 308.290 95.105 ;
        RECT 306.605 94.905 306.925 94.965 ;
        RECT 308.000 94.920 308.290 94.965 ;
        RECT 302.940 94.765 303.230 94.810 ;
        RECT 285.445 94.625 293.955 94.765 ;
        RECT 285.445 94.565 285.765 94.625 ;
        RECT 277.640 94.240 277.930 94.470 ;
        RECT 278.545 94.225 278.865 94.485 ;
        RECT 281.780 94.425 282.070 94.470 ;
        RECT 282.685 94.425 283.005 94.485 ;
        RECT 279.095 94.285 283.005 94.425 ;
        RECT 254.625 94.085 254.945 94.145 ;
        RECT 250.575 93.945 254.945 94.085 ;
        RECT 248.645 93.885 248.965 93.945 ;
        RECT 254.625 93.885 254.945 93.945 ;
        RECT 257.845 94.085 258.165 94.145 ;
        RECT 265.205 94.085 265.525 94.145 ;
        RECT 257.845 93.945 265.525 94.085 ;
        RECT 277.255 94.085 277.395 94.225 ;
        RECT 279.095 94.085 279.235 94.285 ;
        RECT 281.780 94.240 282.070 94.285 ;
        RECT 282.685 94.225 283.005 94.285 ;
        RECT 283.145 94.225 283.465 94.485 ;
        RECT 293.265 94.225 293.585 94.485 ;
        RECT 293.815 94.425 293.955 94.625 ;
        RECT 295.565 94.625 300.855 94.765 ;
        RECT 301.175 94.625 303.230 94.765 ;
        RECT 295.565 94.565 295.885 94.625 ;
        RECT 298.800 94.425 299.090 94.470 ;
        RECT 301.175 94.425 301.315 94.625 ;
        RECT 302.940 94.580 303.230 94.625 ;
        RECT 303.385 94.765 303.705 94.825 ;
        RECT 303.385 94.625 307.295 94.765 ;
        RECT 303.385 94.565 303.705 94.625 ;
        RECT 293.815 94.285 301.315 94.425 ;
        RECT 298.800 94.240 299.090 94.285 ;
        RECT 302.465 94.225 302.785 94.485 ;
        RECT 304.780 94.425 305.070 94.470 ;
        RECT 305.685 94.425 306.005 94.485 ;
        RECT 307.155 94.470 307.295 94.625 ;
        RECT 304.780 94.285 306.005 94.425 ;
        RECT 304.780 94.240 305.070 94.285 ;
        RECT 305.685 94.225 306.005 94.285 ;
        RECT 307.080 94.240 307.370 94.470 ;
        RECT 287.745 94.085 288.065 94.145 ;
        RECT 277.255 93.945 279.235 94.085 ;
        RECT 283.695 93.945 288.065 94.085 ;
        RECT 257.845 93.885 258.165 93.945 ;
        RECT 265.205 93.885 265.525 93.945 ;
        RECT 247.265 93.745 247.585 93.805 ;
        RECT 273.485 93.745 273.805 93.805 ;
        RECT 283.695 93.745 283.835 93.945 ;
        RECT 287.745 93.885 288.065 93.945 ;
        RECT 294.660 93.900 294.950 94.130 ;
        RECT 247.265 93.605 273.805 93.745 ;
        RECT 247.265 93.545 247.585 93.605 ;
        RECT 273.485 93.545 273.805 93.605 ;
        RECT 274.035 93.605 283.835 93.745 ;
        RECT 284.080 93.745 284.370 93.790 ;
        RECT 294.735 93.745 294.875 93.900 ;
        RECT 299.705 93.885 300.025 94.145 ;
        RECT 303.400 93.900 303.690 94.130 ;
        RECT 299.795 93.745 299.935 93.885 ;
        RECT 303.475 93.745 303.615 93.900 ;
        RECT 284.080 93.605 299.935 93.745 ;
        RECT 303.015 93.605 303.615 93.745 ;
        RECT 248.185 93.405 248.505 93.465 ;
        RECT 246.895 93.265 248.505 93.405 ;
        RECT 241.745 93.205 242.065 93.265 ;
        RECT 245.885 93.205 246.205 93.265 ;
        RECT 248.185 93.205 248.505 93.265 ;
        RECT 250.485 93.205 250.805 93.465 ;
        RECT 250.945 93.405 251.265 93.465 ;
        RECT 274.035 93.405 274.175 93.605 ;
        RECT 284.080 93.560 284.370 93.605 ;
        RECT 250.945 93.265 274.175 93.405 ;
        RECT 274.405 93.405 274.725 93.465 ;
        RECT 282.240 93.405 282.530 93.450 ;
        RECT 274.405 93.265 282.530 93.405 ;
        RECT 250.945 93.205 251.265 93.265 ;
        RECT 274.405 93.205 274.725 93.265 ;
        RECT 282.240 93.220 282.530 93.265 ;
        RECT 291.440 93.405 291.730 93.450 ;
        RECT 293.725 93.405 294.045 93.465 ;
        RECT 291.440 93.265 294.045 93.405 ;
        RECT 291.440 93.220 291.730 93.265 ;
        RECT 293.725 93.205 294.045 93.265 ;
        RECT 298.325 93.405 298.645 93.465 ;
        RECT 303.015 93.405 303.155 93.605 ;
        RECT 298.325 93.265 303.155 93.405 ;
        RECT 298.325 93.205 298.645 93.265 ;
        RECT 162.095 92.585 311.135 93.065 ;
        RECT 193.445 92.385 193.765 92.445 ;
        RECT 215.065 92.385 215.385 92.445 ;
        RECT 182.495 92.245 193.765 92.385 ;
        RECT 165.385 92.045 165.705 92.105 ;
        RECT 182.495 92.045 182.635 92.245 ;
        RECT 193.445 92.185 193.765 92.245 ;
        RECT 196.295 92.245 215.385 92.385 ;
        RECT 165.385 91.905 182.635 92.045 ;
        RECT 165.385 91.845 165.705 91.905 ;
        RECT 172.285 91.705 172.605 91.765 ;
        RECT 182.495 91.750 182.635 91.905 ;
        RECT 184.210 92.045 184.500 92.090 ;
        RECT 186.100 92.045 186.390 92.090 ;
        RECT 189.220 92.045 189.510 92.090 ;
        RECT 184.210 91.905 189.510 92.045 ;
        RECT 184.210 91.860 184.500 91.905 ;
        RECT 186.100 91.860 186.390 91.905 ;
        RECT 189.220 91.860 189.510 91.905 ;
        RECT 174.140 91.705 174.430 91.750 ;
        RECT 178.280 91.705 178.570 91.750 ;
        RECT 172.285 91.565 178.570 91.705 ;
        RECT 172.285 91.505 172.605 91.565 ;
        RECT 174.140 91.520 174.430 91.565 ;
        RECT 178.280 91.520 178.570 91.565 ;
        RECT 182.420 91.520 182.710 91.750 ;
        RECT 184.720 91.705 185.010 91.750 ;
        RECT 187.925 91.705 188.245 91.765 ;
        RECT 184.720 91.565 188.245 91.705 ;
        RECT 184.720 91.520 185.010 91.565 ;
        RECT 187.925 91.505 188.245 91.565 ;
        RECT 192.065 91.505 192.385 91.765 ;
        RECT 173.220 91.365 173.510 91.410 ;
        RECT 174.585 91.365 174.905 91.425 ;
        RECT 173.220 91.225 183.095 91.365 ;
        RECT 173.220 91.180 173.510 91.225 ;
        RECT 174.585 91.165 174.905 91.225 ;
        RECT 172.760 91.025 173.050 91.070 ;
        RECT 176.885 91.025 177.205 91.085 ;
        RECT 172.760 90.885 177.205 91.025 ;
        RECT 172.760 90.840 173.050 90.885 ;
        RECT 176.885 90.825 177.205 90.885 ;
        RECT 177.360 91.025 177.650 91.070 ;
        RECT 179.660 91.025 179.950 91.070 ;
        RECT 177.360 90.885 179.950 91.025 ;
        RECT 182.955 91.025 183.095 91.225 ;
        RECT 183.325 91.165 183.645 91.425 ;
        RECT 183.805 91.365 184.095 91.410 ;
        RECT 185.640 91.365 185.930 91.410 ;
        RECT 189.220 91.365 189.510 91.410 ;
        RECT 183.805 91.225 189.510 91.365 ;
        RECT 183.805 91.180 184.095 91.225 ;
        RECT 185.640 91.180 185.930 91.225 ;
        RECT 189.220 91.180 189.510 91.225 ;
        RECT 186.085 91.025 186.405 91.085 ;
        RECT 190.300 91.070 190.590 91.385 ;
        RECT 194.840 91.365 195.130 91.410 ;
        RECT 195.285 91.365 195.605 91.425 ;
        RECT 194.840 91.225 195.605 91.365 ;
        RECT 194.840 91.180 195.130 91.225 ;
        RECT 195.285 91.165 195.605 91.225 ;
        RECT 195.745 91.165 196.065 91.425 ;
        RECT 196.295 91.410 196.435 92.245 ;
        RECT 215.065 92.185 215.385 92.245 ;
        RECT 227.025 92.385 227.345 92.445 ;
        RECT 228.865 92.385 229.185 92.445 ;
        RECT 227.025 92.245 229.185 92.385 ;
        RECT 227.025 92.185 227.345 92.245 ;
        RECT 228.865 92.185 229.185 92.245 ;
        RECT 233.005 92.385 233.325 92.445 ;
        RECT 250.945 92.385 251.265 92.445 ;
        RECT 233.005 92.245 251.265 92.385 ;
        RECT 233.005 92.185 233.325 92.245 ;
        RECT 250.945 92.185 251.265 92.245 ;
        RECT 261.985 92.185 262.305 92.445 ;
        RECT 266.125 92.385 266.445 92.445 ;
        RECT 279.925 92.385 280.245 92.445 ;
        RECT 266.125 92.245 280.245 92.385 ;
        RECT 266.125 92.185 266.445 92.245 ;
        RECT 279.925 92.185 280.245 92.245 ;
        RECT 290.505 92.385 290.825 92.445 ;
        RECT 302.940 92.385 303.230 92.430 ;
        RECT 290.505 92.245 303.230 92.385 ;
        RECT 290.505 92.185 290.825 92.245 ;
        RECT 302.940 92.200 303.230 92.245 ;
        RECT 308.905 92.185 309.225 92.445 ;
        RECT 204.485 92.045 204.805 92.105 ;
        RECT 204.960 92.045 205.250 92.090 ;
        RECT 214.605 92.045 214.925 92.105 ;
        RECT 230.705 92.045 231.025 92.105 ;
        RECT 244.980 92.045 245.270 92.090 ;
        RECT 204.485 91.905 214.925 92.045 ;
        RECT 204.485 91.845 204.805 91.905 ;
        RECT 204.960 91.860 205.250 91.905 ;
        RECT 214.605 91.845 214.925 91.905 ;
        RECT 228.495 91.905 230.475 92.045 ;
        RECT 205.865 91.705 206.185 91.765 ;
        RECT 205.865 91.565 210.235 91.705 ;
        RECT 205.865 91.505 206.185 91.565 ;
        RECT 196.220 91.180 196.510 91.410 ;
        RECT 196.680 91.365 196.970 91.410 ;
        RECT 200.345 91.365 200.665 91.425 ;
        RECT 196.680 91.225 200.665 91.365 ;
        RECT 196.680 91.180 196.970 91.225 ;
        RECT 200.345 91.165 200.665 91.225 ;
        RECT 204.040 91.180 204.330 91.410 ;
        RECT 206.340 91.365 206.630 91.410 ;
        RECT 207.245 91.365 207.565 91.425 ;
        RECT 206.340 91.225 207.565 91.365 ;
        RECT 206.340 91.180 206.630 91.225 ;
        RECT 182.955 90.885 186.405 91.025 ;
        RECT 177.360 90.840 177.650 90.885 ;
        RECT 179.660 90.840 179.950 90.885 ;
        RECT 186.085 90.825 186.405 90.885 ;
        RECT 187.000 91.025 187.650 91.070 ;
        RECT 190.300 91.025 190.890 91.070 ;
        RECT 191.145 91.025 191.465 91.085 ;
        RECT 187.000 90.885 191.465 91.025 ;
        RECT 187.000 90.840 187.650 90.885 ;
        RECT 190.600 90.840 190.890 90.885 ;
        RECT 191.145 90.825 191.465 90.885 ;
        RECT 191.605 91.025 191.925 91.085 ;
        RECT 204.115 91.025 204.255 91.180 ;
        RECT 207.245 91.165 207.565 91.225 ;
        RECT 207.720 91.180 208.010 91.410 ;
        RECT 191.605 90.885 204.255 91.025 ;
        RECT 207.795 91.025 207.935 91.180 ;
        RECT 209.085 91.165 209.405 91.425 ;
        RECT 210.095 91.410 210.235 91.565 ;
        RECT 210.465 91.505 210.785 91.765 ;
        RECT 210.020 91.180 210.310 91.410 ;
        RECT 210.925 91.165 211.245 91.425 ;
        RECT 211.385 91.365 211.705 91.425 ;
        RECT 211.860 91.365 212.150 91.410 ;
        RECT 211.385 91.225 212.150 91.365 ;
        RECT 211.385 91.165 211.705 91.225 ;
        RECT 211.860 91.180 212.150 91.225 ;
        RECT 212.780 91.365 213.070 91.410 ;
        RECT 215.985 91.365 216.305 91.425 ;
        RECT 212.780 91.225 216.305 91.365 ;
        RECT 212.780 91.180 213.070 91.225 ;
        RECT 215.985 91.165 216.305 91.225 ;
        RECT 223.345 91.365 223.665 91.425 ;
        RECT 224.280 91.365 224.570 91.410 ;
        RECT 223.345 91.225 224.570 91.365 ;
        RECT 223.345 91.165 223.665 91.225 ;
        RECT 224.280 91.180 224.570 91.225 ;
        RECT 224.725 91.365 225.045 91.425 ;
        RECT 226.120 91.365 226.410 91.410 ;
        RECT 226.565 91.365 226.885 91.425 ;
        RECT 227.945 91.410 228.265 91.425 ;
        RECT 228.495 91.410 228.635 91.905 ;
        RECT 229.325 91.705 229.645 91.765 ;
        RECT 230.335 91.705 230.475 91.905 ;
        RECT 230.705 91.905 245.270 92.045 ;
        RECT 230.705 91.845 231.025 91.905 ;
        RECT 244.980 91.860 245.270 91.905 ;
        RECT 245.425 92.045 245.745 92.105 ;
        RECT 286.380 92.045 286.670 92.090 ;
        RECT 245.425 91.905 286.670 92.045 ;
        RECT 245.425 91.845 245.745 91.905 ;
        RECT 286.380 91.860 286.670 91.905 ;
        RECT 289.240 92.045 289.530 92.090 ;
        RECT 292.360 92.045 292.650 92.090 ;
        RECT 294.250 92.045 294.540 92.090 ;
        RECT 289.240 91.905 294.540 92.045 ;
        RECT 289.240 91.860 289.530 91.905 ;
        RECT 292.360 91.860 292.650 91.905 ;
        RECT 294.250 91.860 294.540 91.905 ;
        RECT 296.485 92.045 296.805 92.105 ;
        RECT 307.065 92.045 307.385 92.105 ;
        RECT 296.485 91.905 307.385 92.045 ;
        RECT 233.005 91.705 233.325 91.765 ;
        RECT 253.705 91.705 254.025 91.765 ;
        RECT 257.845 91.705 258.165 91.765 ;
        RECT 266.125 91.705 266.445 91.765 ;
        RECT 229.325 91.565 229.990 91.705 ;
        RECT 230.335 91.565 233.325 91.705 ;
        RECT 229.325 91.505 229.645 91.565 ;
        RECT 229.850 91.410 229.990 91.565 ;
        RECT 227.935 91.365 228.265 91.410 ;
        RECT 224.725 91.225 225.875 91.365 ;
        RECT 224.725 91.165 225.045 91.225 ;
        RECT 207.795 90.885 221.505 91.025 ;
        RECT 191.605 90.825 191.925 90.885 ;
        RECT 167.225 90.685 167.545 90.745 ;
        RECT 170.920 90.685 171.210 90.730 ;
        RECT 167.225 90.545 171.210 90.685 ;
        RECT 167.225 90.485 167.545 90.545 ;
        RECT 170.920 90.500 171.210 90.545 ;
        RECT 175.045 90.685 175.365 90.745 ;
        RECT 175.520 90.685 175.810 90.730 ;
        RECT 175.045 90.545 175.810 90.685 ;
        RECT 175.045 90.485 175.365 90.545 ;
        RECT 175.520 90.500 175.810 90.545 ;
        RECT 175.965 90.685 176.285 90.745 ;
        RECT 177.820 90.685 178.110 90.730 ;
        RECT 187.925 90.685 188.245 90.745 ;
        RECT 175.965 90.545 188.245 90.685 ;
        RECT 175.965 90.485 176.285 90.545 ;
        RECT 177.820 90.500 178.110 90.545 ;
        RECT 187.925 90.485 188.245 90.545 ;
        RECT 198.045 90.485 198.365 90.745 ;
        RECT 203.565 90.685 203.885 90.745 ;
        RECT 206.800 90.685 207.090 90.730 ;
        RECT 203.565 90.545 207.090 90.685 ;
        RECT 203.565 90.485 203.885 90.545 ;
        RECT 206.800 90.500 207.090 90.545 ;
        RECT 207.705 90.685 208.025 90.745 ;
        RECT 208.640 90.685 208.930 90.730 ;
        RECT 207.705 90.545 208.930 90.685 ;
        RECT 207.705 90.485 208.025 90.545 ;
        RECT 208.640 90.500 208.930 90.545 ;
        RECT 214.605 90.685 214.925 90.745 ;
        RECT 219.205 90.685 219.525 90.745 ;
        RECT 214.605 90.545 219.525 90.685 ;
        RECT 221.365 90.685 221.505 90.885 ;
        RECT 225.185 90.825 225.505 91.085 ;
        RECT 225.735 91.025 225.875 91.225 ;
        RECT 226.120 91.225 226.885 91.365 ;
        RECT 227.750 91.225 228.265 91.365 ;
        RECT 226.120 91.180 226.410 91.225 ;
        RECT 226.565 91.165 226.885 91.225 ;
        RECT 227.935 91.180 228.265 91.225 ;
        RECT 228.420 91.180 228.710 91.410 ;
        RECT 229.795 91.180 230.085 91.410 ;
        RECT 230.260 91.365 230.550 91.410 ;
        RECT 230.705 91.365 231.025 91.425 ;
        RECT 230.260 91.225 231.025 91.365 ;
        RECT 230.260 91.180 230.550 91.225 ;
        RECT 227.945 91.165 228.265 91.180 ;
        RECT 230.705 91.165 231.025 91.225 ;
        RECT 231.625 91.165 231.945 91.425 ;
        RECT 232.175 91.410 232.315 91.565 ;
        RECT 233.005 91.505 233.325 91.565 ;
        RECT 242.755 91.565 247.495 91.705 ;
        RECT 232.100 91.180 232.390 91.410 ;
        RECT 232.545 91.165 232.865 91.425 ;
        RECT 233.480 91.180 233.770 91.410 ;
        RECT 240.825 91.365 241.145 91.425 ;
        RECT 242.755 91.410 242.895 91.565 ;
        RECT 245.885 91.410 246.205 91.425 ;
        RECT 242.220 91.365 242.510 91.410 ;
        RECT 240.825 91.225 242.510 91.365 ;
        RECT 225.735 90.885 228.180 91.025 ;
        RECT 223.360 90.685 223.650 90.730 ;
        RECT 221.365 90.545 223.650 90.685 ;
        RECT 214.605 90.485 214.925 90.545 ;
        RECT 219.205 90.485 219.525 90.545 ;
        RECT 223.360 90.500 223.650 90.545 ;
        RECT 224.265 90.685 224.585 90.745 ;
        RECT 227.040 90.685 227.330 90.730 ;
        RECT 224.265 90.545 227.330 90.685 ;
        RECT 228.040 90.685 228.180 90.885 ;
        RECT 228.865 90.825 229.185 91.085 ;
        RECT 233.555 91.025 233.695 91.180 ;
        RECT 240.825 91.165 241.145 91.225 ;
        RECT 242.220 91.180 242.510 91.225 ;
        RECT 242.680 91.180 242.970 91.410 ;
        RECT 244.520 91.365 244.810 91.410 ;
        RECT 245.875 91.365 246.205 91.410 ;
        RECT 244.520 91.225 245.425 91.365 ;
        RECT 245.690 91.225 246.205 91.365 ;
        RECT 247.355 91.410 247.495 91.565 ;
        RECT 253.705 91.565 258.165 91.705 ;
        RECT 253.705 91.505 254.025 91.565 ;
        RECT 257.845 91.505 258.165 91.565 ;
        RECT 259.775 91.565 266.445 91.705 ;
        RECT 247.725 91.410 248.045 91.425 ;
        RECT 247.355 91.225 248.045 91.410 ;
        RECT 244.520 91.180 244.810 91.225 ;
        RECT 230.335 90.885 233.695 91.025 ;
        RECT 230.335 90.685 230.475 90.885 ;
        RECT 243.125 90.825 243.445 91.085 ;
        RECT 243.585 91.070 243.905 91.085 ;
        RECT 243.585 90.840 244.020 91.070 ;
        RECT 243.585 90.825 243.905 90.840 ;
        RECT 228.040 90.545 230.475 90.685 ;
        RECT 224.265 90.485 224.585 90.545 ;
        RECT 227.040 90.500 227.330 90.545 ;
        RECT 230.705 90.485 231.025 90.745 ;
        RECT 231.165 90.685 231.485 90.745 ;
        RECT 241.300 90.685 241.590 90.730 ;
        RECT 231.165 90.545 241.590 90.685 ;
        RECT 245.285 90.685 245.425 91.225 ;
        RECT 245.875 91.180 246.205 91.225 ;
        RECT 247.460 91.180 248.045 91.225 ;
        RECT 245.885 91.165 246.205 91.180 ;
        RECT 247.725 91.165 248.045 91.180 ;
        RECT 248.185 91.165 248.505 91.425 ;
        RECT 257.385 91.365 257.705 91.425 ;
        RECT 259.775 91.410 259.915 91.565 ;
        RECT 266.125 91.505 266.445 91.565 ;
        RECT 281.765 91.505 282.085 91.765 ;
        RECT 286.455 91.705 286.595 91.860 ;
        RECT 296.485 91.845 296.805 91.905 ;
        RECT 307.065 91.845 307.385 91.905 ;
        RECT 293.265 91.705 293.585 91.765 ;
        RECT 286.455 91.565 293.585 91.705 ;
        RECT 293.265 91.505 293.585 91.565 ;
        RECT 293.725 91.505 294.045 91.765 ;
        RECT 298.340 91.705 298.630 91.750 ;
        RECT 298.785 91.705 299.105 91.765 ;
        RECT 298.340 91.565 299.105 91.705 ;
        RECT 298.340 91.520 298.630 91.565 ;
        RECT 298.785 91.505 299.105 91.565 ;
        RECT 299.260 91.705 299.550 91.750 ;
        RECT 299.705 91.705 300.025 91.765 ;
        RECT 299.260 91.565 300.025 91.705 ;
        RECT 299.260 91.520 299.550 91.565 ;
        RECT 299.705 91.505 300.025 91.565 ;
        RECT 258.780 91.365 259.070 91.410 ;
        RECT 257.385 91.225 259.070 91.365 ;
        RECT 257.385 91.165 257.705 91.225 ;
        RECT 258.780 91.180 259.070 91.225 ;
        RECT 259.520 91.225 259.915 91.410 ;
        RECT 261.065 91.410 261.385 91.425 ;
        RECT 259.520 91.180 259.810 91.225 ;
        RECT 261.065 91.180 261.395 91.410 ;
        RECT 262.460 91.180 262.750 91.410 ;
        RECT 263.840 91.365 264.130 91.410 ;
        RECT 262.995 91.225 264.130 91.365 ;
        RECT 261.065 91.165 261.385 91.180 ;
        RECT 246.360 90.840 246.650 91.070 ;
        RECT 246.820 91.025 247.110 91.070 ;
        RECT 248.645 91.025 248.965 91.085 ;
        RECT 260.145 91.025 260.465 91.085 ;
        RECT 246.820 90.885 260.465 91.025 ;
        RECT 246.820 90.840 247.110 90.885 ;
        RECT 246.435 90.685 246.575 90.840 ;
        RECT 247.815 90.745 247.955 90.885 ;
        RECT 248.645 90.825 248.965 90.885 ;
        RECT 260.145 90.825 260.465 90.885 ;
        RECT 260.620 91.025 260.910 91.070 ;
        RECT 262.535 91.025 262.675 91.180 ;
        RECT 260.620 90.885 262.675 91.025 ;
        RECT 260.620 90.840 260.910 90.885 ;
        RECT 247.265 90.685 247.585 90.745 ;
        RECT 245.285 90.545 247.585 90.685 ;
        RECT 231.165 90.485 231.485 90.545 ;
        RECT 241.300 90.500 241.590 90.545 ;
        RECT 247.265 90.485 247.585 90.545 ;
        RECT 247.725 90.485 248.045 90.745 ;
        RECT 259.685 90.685 260.005 90.745 ;
        RECT 260.695 90.685 260.835 90.840 ;
        RECT 259.685 90.545 260.835 90.685 ;
        RECT 261.065 90.685 261.385 90.745 ;
        RECT 262.995 90.685 263.135 91.225 ;
        RECT 263.840 91.180 264.130 91.225 ;
        RECT 264.300 91.365 264.590 91.410 ;
        RECT 265.205 91.365 265.525 91.425 ;
        RECT 264.300 91.225 265.525 91.365 ;
        RECT 264.300 91.180 264.590 91.225 ;
        RECT 263.380 90.840 263.670 91.070 ;
        RECT 263.915 91.025 264.055 91.180 ;
        RECT 265.205 91.165 265.525 91.225 ;
        RECT 265.680 91.180 265.970 91.410 ;
        RECT 265.755 91.025 265.895 91.180 ;
        RECT 267.505 91.165 267.825 91.425 ;
        RECT 278.085 91.365 278.405 91.425 ;
        RECT 279.480 91.365 279.770 91.410 ;
        RECT 278.085 91.225 279.770 91.365 ;
        RECT 278.085 91.165 278.405 91.225 ;
        RECT 279.480 91.180 279.770 91.225 ;
        RECT 279.925 91.165 280.245 91.425 ;
        RECT 280.845 91.410 281.165 91.425 ;
        RECT 280.845 91.180 281.280 91.410 ;
        RECT 288.205 91.385 288.525 91.425 ;
        RECT 280.845 91.165 281.165 91.180 ;
        RECT 288.160 91.165 288.525 91.385 ;
        RECT 289.240 91.365 289.530 91.410 ;
        RECT 292.820 91.365 293.110 91.410 ;
        RECT 294.655 91.365 294.945 91.410 ;
        RECT 289.240 91.225 294.945 91.365 ;
        RECT 289.240 91.180 289.530 91.225 ;
        RECT 292.820 91.180 293.110 91.225 ;
        RECT 294.655 91.180 294.945 91.225 ;
        RECT 295.105 91.165 295.425 91.425 ;
        RECT 297.865 91.165 298.185 91.425 ;
        RECT 302.020 91.365 302.310 91.410 ;
        RECT 298.875 91.225 302.310 91.365 ;
        RECT 263.915 90.885 265.895 91.025 ;
        RECT 261.065 90.545 263.135 90.685 ;
        RECT 263.455 90.685 263.595 90.840 ;
        RECT 266.585 90.825 266.905 91.085 ;
        RECT 267.045 90.825 267.365 91.085 ;
        RECT 279.005 91.025 279.325 91.085 ;
        RECT 288.160 91.070 288.450 91.165 ;
        RECT 298.875 91.085 299.015 91.225 ;
        RECT 302.020 91.180 302.310 91.225 ;
        RECT 308.000 91.365 308.290 91.410 ;
        RECT 309.825 91.365 310.145 91.425 ;
        RECT 308.000 91.225 310.145 91.365 ;
        RECT 308.000 91.180 308.290 91.225 ;
        RECT 309.825 91.165 310.145 91.225 ;
        RECT 280.400 91.025 280.690 91.070 ;
        RECT 267.595 90.885 279.325 91.025 ;
        RECT 264.745 90.685 265.065 90.745 ;
        RECT 263.455 90.545 265.065 90.685 ;
        RECT 259.685 90.485 260.005 90.545 ;
        RECT 261.065 90.485 261.385 90.545 ;
        RECT 264.745 90.485 265.065 90.545 ;
        RECT 265.220 90.685 265.510 90.730 ;
        RECT 267.595 90.685 267.735 90.885 ;
        RECT 279.005 90.825 279.325 90.885 ;
        RECT 279.555 90.885 280.690 91.025 ;
        RECT 279.555 90.745 279.695 90.885 ;
        RECT 280.400 90.840 280.690 90.885 ;
        RECT 287.860 91.025 288.450 91.070 ;
        RECT 291.100 91.025 291.750 91.070 ;
        RECT 287.860 90.885 291.750 91.025 ;
        RECT 287.860 90.840 288.150 90.885 ;
        RECT 291.100 90.840 291.750 90.885 ;
        RECT 298.785 90.825 299.105 91.085 ;
        RECT 302.465 91.025 302.785 91.085 ;
        RECT 304.780 91.025 305.070 91.070 ;
        RECT 302.465 90.885 305.070 91.025 ;
        RECT 302.465 90.825 302.785 90.885 ;
        RECT 304.780 90.840 305.070 90.885 ;
        RECT 265.220 90.545 267.735 90.685 ;
        RECT 268.440 90.685 268.730 90.730 ;
        RECT 268.885 90.685 269.205 90.745 ;
        RECT 268.440 90.545 269.205 90.685 ;
        RECT 265.220 90.500 265.510 90.545 ;
        RECT 268.440 90.500 268.730 90.545 ;
        RECT 268.885 90.485 269.205 90.545 ;
        RECT 278.545 90.485 278.865 90.745 ;
        RECT 279.465 90.485 279.785 90.745 ;
        RECT 296.040 90.685 296.330 90.730 ;
        RECT 296.485 90.685 296.805 90.745 ;
        RECT 296.040 90.545 296.805 90.685 ;
        RECT 296.040 90.500 296.330 90.545 ;
        RECT 296.485 90.485 296.805 90.545 ;
        RECT 300.165 90.685 300.485 90.745 ;
        RECT 305.240 90.685 305.530 90.730 ;
        RECT 300.165 90.545 305.530 90.685 ;
        RECT 300.165 90.485 300.485 90.545 ;
        RECT 305.240 90.500 305.530 90.545 ;
        RECT 162.095 89.865 311.135 90.345 ;
        RECT 165.845 89.665 166.165 89.725 ;
        RECT 180.565 89.665 180.885 89.725 ;
        RECT 183.325 89.665 183.645 89.725 ;
        RECT 165.845 89.525 183.645 89.665 ;
        RECT 165.845 89.465 166.165 89.525 ;
        RECT 169.180 89.325 169.470 89.370 ;
        RECT 171.825 89.325 172.145 89.385 ;
        RECT 172.420 89.325 173.070 89.370 ;
        RECT 169.180 89.185 173.070 89.325 ;
        RECT 169.180 89.140 169.770 89.185 ;
        RECT 169.480 88.825 169.770 89.140 ;
        RECT 171.825 89.125 172.145 89.185 ;
        RECT 172.420 89.140 173.070 89.185 ;
        RECT 175.045 89.125 175.365 89.385 ;
        RECT 176.515 89.030 176.655 89.525 ;
        RECT 180.565 89.465 180.885 89.525 ;
        RECT 183.325 89.465 183.645 89.525 ;
        RECT 193.000 89.665 193.290 89.710 ;
        RECT 195.745 89.665 196.065 89.725 ;
        RECT 210.925 89.665 211.245 89.725 ;
        RECT 227.025 89.665 227.345 89.725 ;
        RECT 193.000 89.525 196.065 89.665 ;
        RECT 193.000 89.480 193.290 89.525 ;
        RECT 195.745 89.465 196.065 89.525 ;
        RECT 200.895 89.525 211.245 89.665 ;
        RECT 176.885 89.325 177.205 89.385 ;
        RECT 181.040 89.325 181.330 89.370 ;
        RECT 189.305 89.325 189.625 89.385 ;
        RECT 191.145 89.325 191.465 89.385 ;
        RECT 176.885 89.185 181.330 89.325 ;
        RECT 176.885 89.125 177.205 89.185 ;
        RECT 181.040 89.140 181.330 89.185 ;
        RECT 185.715 89.185 191.465 89.325 ;
        RECT 170.560 88.985 170.850 89.030 ;
        RECT 174.140 88.985 174.430 89.030 ;
        RECT 175.975 88.985 176.265 89.030 ;
        RECT 170.560 88.845 176.265 88.985 ;
        RECT 170.560 88.800 170.850 88.845 ;
        RECT 174.140 88.800 174.430 88.845 ;
        RECT 175.975 88.800 176.265 88.845 ;
        RECT 176.440 88.800 176.730 89.030 ;
        RECT 177.345 88.985 177.665 89.045 ;
        RECT 178.740 88.985 179.030 89.030 ;
        RECT 179.645 88.985 179.965 89.045 ;
        RECT 185.715 89.030 185.855 89.185 ;
        RECT 189.305 89.125 189.625 89.185 ;
        RECT 191.145 89.125 191.465 89.185 ;
        RECT 193.445 89.325 193.765 89.385 ;
        RECT 193.920 89.325 194.210 89.370 ;
        RECT 193.445 89.185 194.210 89.325 ;
        RECT 193.445 89.125 193.765 89.185 ;
        RECT 193.920 89.140 194.210 89.185 ;
        RECT 184.720 88.985 185.010 89.030 ;
        RECT 177.345 88.845 179.965 88.985 ;
        RECT 177.345 88.785 177.665 88.845 ;
        RECT 178.740 88.800 179.030 88.845 ;
        RECT 179.645 88.785 179.965 88.845 ;
        RECT 180.195 88.845 185.010 88.985 ;
        RECT 165.385 88.645 165.705 88.705 ;
        RECT 167.700 88.645 167.990 88.690 ;
        RECT 165.385 88.505 167.990 88.645 ;
        RECT 165.385 88.445 165.705 88.505 ;
        RECT 167.700 88.460 167.990 88.505 ;
        RECT 172.285 88.645 172.605 88.705 ;
        RECT 172.285 88.505 178.955 88.645 ;
        RECT 172.285 88.445 172.605 88.505 ;
        RECT 170.560 88.305 170.850 88.350 ;
        RECT 173.680 88.305 173.970 88.350 ;
        RECT 175.570 88.305 175.860 88.350 ;
        RECT 178.815 88.305 178.955 88.505 ;
        RECT 179.185 88.445 179.505 88.705 ;
        RECT 180.195 88.690 180.335 88.845 ;
        RECT 184.720 88.800 185.010 88.845 ;
        RECT 185.640 88.800 185.930 89.030 ;
        RECT 186.545 88.985 186.865 89.045 ;
        RECT 191.605 88.985 191.925 89.045 ;
        RECT 186.545 88.845 191.925 88.985 ;
        RECT 186.545 88.785 186.865 88.845 ;
        RECT 191.605 88.785 191.925 88.845 ;
        RECT 194.840 88.985 195.130 89.030 ;
        RECT 195.745 88.985 196.065 89.045 ;
        RECT 200.895 89.030 201.035 89.525 ;
        RECT 210.925 89.465 211.245 89.525 ;
        RECT 226.195 89.525 227.345 89.665 ;
        RECT 202.660 89.325 202.950 89.370 ;
        RECT 224.265 89.325 224.585 89.385 ;
        RECT 202.660 89.185 207.015 89.325 ;
        RECT 202.660 89.140 202.950 89.185 ;
        RECT 200.820 88.985 201.110 89.030 ;
        RECT 194.840 88.845 201.110 88.985 ;
        RECT 194.840 88.800 195.130 88.845 ;
        RECT 195.745 88.785 196.065 88.845 ;
        RECT 200.820 88.800 201.110 88.845 ;
        RECT 201.725 88.785 202.045 89.045 ;
        RECT 203.105 88.785 203.425 89.045 ;
        RECT 203.565 88.785 203.885 89.045 ;
        RECT 204.485 88.785 204.805 89.045 ;
        RECT 206.875 89.030 207.015 89.185 ;
        RECT 207.335 89.185 224.585 89.325 ;
        RECT 207.335 89.030 207.475 89.185 ;
        RECT 224.265 89.125 224.585 89.185 ;
        RECT 205.880 88.985 206.170 89.030 ;
        RECT 205.880 88.845 206.280 88.985 ;
        RECT 205.880 88.800 206.170 88.845 ;
        RECT 206.800 88.800 207.090 89.030 ;
        RECT 207.260 88.800 207.550 89.030 ;
        RECT 180.120 88.460 180.410 88.690 ;
        RECT 183.800 88.645 184.090 88.690 ;
        RECT 183.415 88.505 184.090 88.645 ;
        RECT 180.195 88.305 180.335 88.460 ;
        RECT 170.560 88.165 175.860 88.305 ;
        RECT 170.560 88.120 170.850 88.165 ;
        RECT 173.680 88.120 173.970 88.165 ;
        RECT 175.570 88.120 175.860 88.165 ;
        RECT 176.515 88.165 178.495 88.305 ;
        RECT 178.815 88.165 180.335 88.305 ;
        RECT 183.415 88.305 183.555 88.505 ;
        RECT 183.800 88.460 184.090 88.505 ;
        RECT 187.005 88.445 187.325 88.705 ;
        RECT 195.285 88.645 195.605 88.705 ;
        RECT 205.955 88.645 206.095 88.800 ;
        RECT 207.705 88.785 208.025 89.045 ;
        RECT 214.145 88.785 214.465 89.045 ;
        RECT 214.605 88.785 214.925 89.045 ;
        RECT 215.540 88.800 215.830 89.030 ;
        RECT 216.000 88.985 216.290 89.030 ;
        RECT 216.905 88.985 217.225 89.045 ;
        RECT 225.645 88.985 225.965 89.045 ;
        RECT 226.195 89.030 226.335 89.525 ;
        RECT 227.025 89.465 227.345 89.525 ;
        RECT 228.880 89.480 229.170 89.710 ;
        RECT 229.785 89.665 230.105 89.725 ;
        RECT 261.065 89.665 261.385 89.725 ;
        RECT 229.785 89.525 261.385 89.665 ;
        RECT 226.565 89.325 226.885 89.385 ;
        RECT 226.565 89.185 227.715 89.325 ;
        RECT 226.565 89.125 226.885 89.185 ;
        RECT 227.575 89.030 227.715 89.185 ;
        RECT 216.000 88.845 217.225 88.985 ;
        RECT 216.000 88.800 216.290 88.845 ;
        RECT 209.085 88.645 209.405 88.705 ;
        RECT 195.285 88.505 209.405 88.645 ;
        RECT 215.615 88.645 215.755 88.800 ;
        RECT 216.905 88.785 217.225 88.845 ;
        RECT 218.835 88.845 225.965 88.985 ;
        RECT 218.835 88.645 218.975 88.845 ;
        RECT 225.645 88.785 225.965 88.845 ;
        RECT 226.120 88.800 226.410 89.030 ;
        RECT 227.040 88.800 227.330 89.030 ;
        RECT 227.500 88.800 227.790 89.030 ;
        RECT 215.615 88.505 218.975 88.645 ;
        RECT 219.205 88.645 219.525 88.705 ;
        RECT 224.725 88.645 225.045 88.705 ;
        RECT 219.205 88.505 225.045 88.645 ;
        RECT 195.285 88.445 195.605 88.505 ;
        RECT 209.085 88.445 209.405 88.505 ;
        RECT 219.205 88.445 219.525 88.505 ;
        RECT 224.725 88.445 225.045 88.505 ;
        RECT 226.565 88.645 226.885 88.705 ;
        RECT 227.115 88.645 227.255 88.800 ;
        RECT 226.565 88.505 227.255 88.645 ;
        RECT 227.575 88.645 227.715 88.800 ;
        RECT 227.945 88.785 228.265 89.045 ;
        RECT 228.955 88.985 229.095 89.480 ;
        RECT 229.785 89.465 230.105 89.525 ;
        RECT 261.065 89.465 261.385 89.525 ;
        RECT 261.525 89.665 261.845 89.725 ;
        RECT 268.440 89.665 268.730 89.710 ;
        RECT 293.265 89.665 293.585 89.725 ;
        RECT 261.525 89.525 266.815 89.665 ;
        RECT 261.525 89.465 261.845 89.525 ;
        RECT 258.305 89.325 258.625 89.385 ;
        RECT 244.595 89.185 258.625 89.325 ;
        RECT 230.260 88.985 230.550 89.030 ;
        RECT 228.955 88.845 230.550 88.985 ;
        RECT 230.260 88.800 230.550 88.845 ;
        RECT 231.165 88.785 231.485 89.045 ;
        RECT 244.595 89.030 244.735 89.185 ;
        RECT 258.305 89.125 258.625 89.185 ;
        RECT 259.685 89.325 260.005 89.385 ;
        RECT 266.675 89.370 266.815 89.525 ;
        RECT 268.440 89.525 278.315 89.665 ;
        RECT 268.440 89.480 268.730 89.525 ;
        RECT 262.460 89.325 262.750 89.370 ;
        RECT 259.685 89.185 262.750 89.325 ;
        RECT 259.685 89.125 260.005 89.185 ;
        RECT 262.460 89.140 262.750 89.185 ;
        RECT 262.995 89.185 265.895 89.325 ;
        RECT 262.995 89.045 263.135 89.185 ;
        RECT 244.520 88.800 244.810 89.030 ;
        RECT 244.965 88.785 245.285 89.045 ;
        RECT 245.900 88.800 246.190 89.030 ;
        RECT 245.425 88.645 245.745 88.705 ;
        RECT 227.575 88.505 245.745 88.645 ;
        RECT 245.975 88.645 246.115 88.800 ;
        RECT 246.345 88.785 246.665 89.045 ;
        RECT 250.485 88.985 250.805 89.045 ;
        RECT 261.080 88.985 261.370 89.030 ;
        RECT 250.485 88.845 261.370 88.985 ;
        RECT 250.485 88.785 250.805 88.845 ;
        RECT 261.080 88.800 261.370 88.845 ;
        RECT 261.820 88.985 262.110 89.030 ;
        RECT 261.820 88.800 262.215 88.985 ;
        RECT 246.805 88.645 247.125 88.705 ;
        RECT 259.225 88.645 259.545 88.705 ;
        RECT 245.975 88.505 259.545 88.645 ;
        RECT 226.565 88.445 226.885 88.505 ;
        RECT 245.425 88.445 245.745 88.505 ;
        RECT 246.805 88.445 247.125 88.505 ;
        RECT 259.225 88.445 259.545 88.505 ;
        RECT 201.725 88.305 202.045 88.365 ;
        RECT 183.415 88.165 202.045 88.305 ;
        RECT 174.125 87.965 174.445 88.025 ;
        RECT 176.515 87.965 176.655 88.165 ;
        RECT 174.125 87.825 176.655 87.965 ;
        RECT 174.125 87.765 174.445 87.825 ;
        RECT 176.885 87.765 177.205 88.025 ;
        RECT 178.355 87.965 178.495 88.165 ;
        RECT 183.415 87.965 183.555 88.165 ;
        RECT 201.725 88.105 202.045 88.165 ;
        RECT 210.005 88.305 210.325 88.365 ;
        RECT 229.340 88.305 229.630 88.350 ;
        RECT 252.785 88.305 253.105 88.365 ;
        RECT 210.005 88.165 229.630 88.305 ;
        RECT 210.005 88.105 210.325 88.165 ;
        RECT 229.340 88.120 229.630 88.165 ;
        RECT 230.335 88.165 253.105 88.305 ;
        RECT 262.075 88.305 262.215 88.800 ;
        RECT 262.905 88.785 263.225 89.045 ;
        RECT 263.610 88.985 263.900 89.030 ;
        RECT 265.205 88.985 265.525 89.045 ;
        RECT 265.755 89.030 265.895 89.185 ;
        RECT 266.600 89.140 266.890 89.370 ;
        RECT 271.185 89.325 271.505 89.385 ;
        RECT 274.405 89.325 274.725 89.385 ;
        RECT 278.175 89.370 278.315 89.525 ;
        RECT 293.265 89.525 306.375 89.665 ;
        RECT 293.265 89.465 293.585 89.525 ;
        RECT 267.595 89.185 274.725 89.325 ;
        RECT 263.610 88.845 265.525 88.985 ;
        RECT 263.610 88.800 263.900 88.845 ;
        RECT 265.205 88.785 265.525 88.845 ;
        RECT 265.680 88.800 265.970 89.030 ;
        RECT 267.045 88.785 267.365 89.045 ;
        RECT 267.595 89.030 267.735 89.185 ;
        RECT 271.185 89.125 271.505 89.185 ;
        RECT 274.405 89.125 274.725 89.185 ;
        RECT 278.100 89.140 278.390 89.370 ;
        RECT 296.485 89.125 296.805 89.385 ;
        RECT 298.780 89.325 299.430 89.370 ;
        RECT 300.165 89.325 300.485 89.385 ;
        RECT 302.380 89.325 302.670 89.370 ;
        RECT 298.780 89.185 302.670 89.325 ;
        RECT 298.780 89.140 299.430 89.185 ;
        RECT 300.165 89.125 300.485 89.185 ;
        RECT 302.080 89.140 302.670 89.185 ;
        RECT 267.520 88.800 267.810 89.030 ;
        RECT 268.885 88.785 269.205 89.045 ;
        RECT 279.005 88.785 279.325 89.045 ;
        RECT 279.480 88.985 279.770 89.030 ;
        RECT 286.825 88.985 287.145 89.045 ;
        RECT 279.480 88.845 287.145 88.985 ;
        RECT 279.480 88.800 279.770 88.845 ;
        RECT 286.825 88.785 287.145 88.845 ;
        RECT 295.585 88.985 295.875 89.030 ;
        RECT 297.420 88.985 297.710 89.030 ;
        RECT 301.000 88.985 301.290 89.030 ;
        RECT 295.585 88.845 301.290 88.985 ;
        RECT 295.585 88.800 295.875 88.845 ;
        RECT 297.420 88.800 297.710 88.845 ;
        RECT 301.000 88.800 301.290 88.845 ;
        RECT 302.080 88.825 302.370 89.140 ;
        RECT 306.235 89.030 306.375 89.525 ;
        RECT 307.065 89.465 307.385 89.725 ;
        RECT 308.920 89.665 309.210 89.710 ;
        RECT 309.365 89.665 309.685 89.725 ;
        RECT 308.920 89.525 309.685 89.665 ;
        RECT 308.920 89.480 309.210 89.525 ;
        RECT 309.365 89.465 309.685 89.525 ;
        RECT 306.160 88.800 306.450 89.030 ;
        RECT 307.985 88.785 308.305 89.045 ;
        RECT 269.360 88.645 269.650 88.690 ;
        RECT 264.375 88.505 269.650 88.645 ;
        RECT 263.825 88.305 264.145 88.365 ;
        RECT 264.375 88.350 264.515 88.505 ;
        RECT 269.360 88.460 269.650 88.505 ;
        RECT 294.645 88.645 294.965 88.705 ;
        RECT 295.120 88.645 295.410 88.690 ;
        RECT 294.645 88.505 295.410 88.645 ;
        RECT 294.645 88.445 294.965 88.505 ;
        RECT 295.120 88.460 295.410 88.505 ;
        RECT 298.325 88.645 298.645 88.705 ;
        RECT 303.845 88.645 304.165 88.705 ;
        RECT 298.325 88.505 304.165 88.645 ;
        RECT 298.325 88.445 298.645 88.505 ;
        RECT 303.845 88.445 304.165 88.505 ;
        RECT 262.075 88.165 264.145 88.305 ;
        RECT 178.355 87.825 183.555 87.965 ;
        RECT 187.925 87.965 188.245 88.025 ;
        RECT 199.885 87.965 200.205 88.025 ;
        RECT 187.925 87.825 200.205 87.965 ;
        RECT 187.925 87.765 188.245 87.825 ;
        RECT 199.885 87.765 200.205 87.825 ;
        RECT 205.420 87.965 205.710 88.010 ;
        RECT 205.865 87.965 206.185 88.025 ;
        RECT 205.420 87.825 206.185 87.965 ;
        RECT 205.420 87.780 205.710 87.825 ;
        RECT 205.865 87.765 206.185 87.825 ;
        RECT 209.085 87.765 209.405 88.025 ;
        RECT 212.765 87.965 213.085 88.025 ;
        RECT 216.920 87.965 217.210 88.010 ;
        RECT 212.765 87.825 217.210 87.965 ;
        RECT 212.765 87.765 213.085 87.825 ;
        RECT 216.920 87.780 217.210 87.825 ;
        RECT 225.645 87.965 225.965 88.025 ;
        RECT 230.335 87.965 230.475 88.165 ;
        RECT 252.785 88.105 253.105 88.165 ;
        RECT 263.825 88.105 264.145 88.165 ;
        RECT 264.300 88.120 264.590 88.350 ;
        RECT 267.045 88.305 267.365 88.365 ;
        RECT 295.990 88.305 296.280 88.350 ;
        RECT 297.880 88.305 298.170 88.350 ;
        RECT 301.000 88.305 301.290 88.350 ;
        RECT 267.045 88.165 281.205 88.305 ;
        RECT 267.045 88.105 267.365 88.165 ;
        RECT 225.645 87.825 230.475 87.965 ;
        RECT 225.645 87.765 225.965 87.825 ;
        RECT 230.705 87.765 231.025 88.025 ;
        RECT 243.585 87.765 243.905 88.025 ;
        RECT 247.265 87.965 247.585 88.025 ;
        RECT 251.405 87.965 251.725 88.025 ;
        RECT 259.685 87.965 260.005 88.025 ;
        RECT 247.265 87.825 260.005 87.965 ;
        RECT 247.265 87.765 247.585 87.825 ;
        RECT 251.405 87.765 251.725 87.825 ;
        RECT 259.685 87.765 260.005 87.825 ;
        RECT 261.985 87.965 262.305 88.025 ;
        RECT 268.900 87.965 269.190 88.010 ;
        RECT 261.985 87.825 269.190 87.965 ;
        RECT 261.985 87.765 262.305 87.825 ;
        RECT 268.900 87.780 269.190 87.825 ;
        RECT 270.725 87.765 271.045 88.025 ;
        RECT 278.545 87.765 278.865 88.025 ;
        RECT 280.385 87.765 280.705 88.025 ;
        RECT 281.065 87.965 281.205 88.165 ;
        RECT 295.990 88.165 301.290 88.305 ;
        RECT 295.990 88.120 296.280 88.165 ;
        RECT 297.880 88.120 298.170 88.165 ;
        RECT 301.000 88.120 301.290 88.165 ;
        RECT 302.005 87.965 302.325 88.025 ;
        RECT 281.065 87.825 302.325 87.965 ;
        RECT 302.005 87.765 302.325 87.825 ;
        RECT 162.095 87.145 311.135 87.625 ;
        RECT 174.125 86.945 174.445 87.005 ;
        RECT 174.600 86.945 174.890 86.990 ;
        RECT 174.125 86.805 174.890 86.945 ;
        RECT 174.125 86.745 174.445 86.805 ;
        RECT 174.600 86.760 174.890 86.805 ;
        RECT 179.645 86.945 179.965 87.005 ;
        RECT 184.260 86.945 184.550 86.990 ;
        RECT 208.625 86.945 208.945 87.005 ;
        RECT 211.385 86.945 211.705 87.005 ;
        RECT 179.645 86.805 211.705 86.945 ;
        RECT 179.645 86.745 179.965 86.805 ;
        RECT 184.260 86.760 184.550 86.805 ;
        RECT 208.625 86.745 208.945 86.805 ;
        RECT 211.385 86.745 211.705 86.805 ;
        RECT 223.805 86.945 224.125 87.005 ;
        RECT 225.645 86.945 225.965 87.005 ;
        RECT 226.565 86.945 226.885 87.005 ;
        RECT 223.805 86.805 226.885 86.945 ;
        RECT 223.805 86.745 224.125 86.805 ;
        RECT 225.645 86.745 225.965 86.805 ;
        RECT 226.565 86.745 226.885 86.805 ;
        RECT 227.945 86.945 228.265 87.005 ;
        RECT 228.865 86.945 229.185 87.005 ;
        RECT 240.365 86.945 240.685 87.005 ;
        RECT 227.945 86.805 240.685 86.945 ;
        RECT 227.945 86.745 228.265 86.805 ;
        RECT 228.865 86.745 229.185 86.805 ;
        RECT 240.365 86.745 240.685 86.805 ;
        RECT 242.665 86.945 242.985 87.005 ;
        RECT 242.665 86.805 249.310 86.945 ;
        RECT 242.665 86.745 242.985 86.805 ;
        RECT 166.730 86.605 167.020 86.650 ;
        RECT 168.620 86.605 168.910 86.650 ;
        RECT 171.740 86.605 172.030 86.650 ;
        RECT 166.730 86.465 172.030 86.605 ;
        RECT 166.730 86.420 167.020 86.465 ;
        RECT 168.620 86.420 168.910 86.465 ;
        RECT 171.740 86.420 172.030 86.465 ;
        RECT 176.390 86.605 176.680 86.650 ;
        RECT 178.280 86.605 178.570 86.650 ;
        RECT 181.400 86.605 181.690 86.650 ;
        RECT 176.390 86.465 181.690 86.605 ;
        RECT 176.390 86.420 176.680 86.465 ;
        RECT 178.280 86.420 178.570 86.465 ;
        RECT 181.400 86.420 181.690 86.465 ;
        RECT 185.165 86.405 185.485 86.665 ;
        RECT 187.925 86.405 188.245 86.665 ;
        RECT 194.825 86.605 195.145 86.665 ;
        RECT 194.825 86.465 210.695 86.605 ;
        RECT 194.825 86.405 195.145 86.465 ;
        RECT 165.845 86.065 166.165 86.325 ;
        RECT 167.225 86.065 167.545 86.325 ;
        RECT 167.685 86.265 168.005 86.325 ;
        RECT 175.520 86.265 175.810 86.310 ;
        RECT 188.385 86.265 188.705 86.325 ;
        RECT 192.985 86.265 193.305 86.325 ;
        RECT 167.685 86.125 193.305 86.265 ;
        RECT 167.685 86.065 168.005 86.125 ;
        RECT 175.520 86.080 175.810 86.125 ;
        RECT 188.385 86.065 188.705 86.125 ;
        RECT 192.985 86.065 193.305 86.125 ;
        RECT 194.455 86.125 201.495 86.265 ;
        RECT 166.325 85.925 166.615 85.970 ;
        RECT 168.160 85.925 168.450 85.970 ;
        RECT 171.740 85.925 172.030 85.970 ;
        RECT 166.325 85.785 172.030 85.925 ;
        RECT 166.325 85.740 166.615 85.785 ;
        RECT 168.160 85.740 168.450 85.785 ;
        RECT 171.740 85.740 172.030 85.785 ;
        RECT 172.820 85.630 173.110 85.945 ;
        RECT 175.985 85.925 176.275 85.970 ;
        RECT 177.820 85.925 178.110 85.970 ;
        RECT 181.400 85.925 181.690 85.970 ;
        RECT 175.985 85.785 181.690 85.925 ;
        RECT 175.985 85.740 176.275 85.785 ;
        RECT 177.820 85.740 178.110 85.785 ;
        RECT 181.400 85.740 181.690 85.785 ;
        RECT 169.520 85.585 170.170 85.630 ;
        RECT 172.820 85.585 173.410 85.630 ;
        RECT 169.520 85.445 175.275 85.585 ;
        RECT 169.520 85.400 170.170 85.445 ;
        RECT 173.120 85.400 173.410 85.445 ;
        RECT 171.825 85.245 172.145 85.305 ;
        RECT 173.755 85.245 173.895 85.445 ;
        RECT 171.825 85.105 173.895 85.245 ;
        RECT 175.135 85.245 175.275 85.445 ;
        RECT 176.885 85.385 177.205 85.645 ;
        RECT 182.480 85.630 182.770 85.945 ;
        RECT 186.100 85.740 186.390 85.970 ;
        RECT 179.180 85.585 179.830 85.630 ;
        RECT 182.480 85.585 183.070 85.630 ;
        RECT 177.435 85.445 183.070 85.585 ;
        RECT 186.175 85.585 186.315 85.740 ;
        RECT 187.005 85.725 187.325 85.985 ;
        RECT 188.860 85.925 189.150 85.970 ;
        RECT 189.305 85.925 189.625 85.985 ;
        RECT 188.860 85.785 189.625 85.925 ;
        RECT 188.860 85.740 189.150 85.785 ;
        RECT 188.935 85.585 189.075 85.740 ;
        RECT 189.305 85.725 189.625 85.785 ;
        RECT 189.780 85.740 190.070 85.970 ;
        RECT 189.855 85.585 189.995 85.740 ;
        RECT 193.445 85.725 193.765 85.985 ;
        RECT 194.455 85.970 194.595 86.125 ;
        RECT 194.380 85.740 194.670 85.970 ;
        RECT 194.825 85.725 195.145 85.985 ;
        RECT 195.760 85.740 196.050 85.970 ;
        RECT 186.175 85.445 189.075 85.585 ;
        RECT 189.395 85.445 189.995 85.585 ;
        RECT 177.435 85.245 177.575 85.445 ;
        RECT 179.180 85.400 179.830 85.445 ;
        RECT 182.780 85.400 183.070 85.445 ;
        RECT 189.395 85.305 189.535 85.445 ;
        RECT 175.135 85.105 177.575 85.245 ;
        RECT 171.825 85.045 172.145 85.105 ;
        RECT 189.305 85.045 189.625 85.305 ;
        RECT 192.540 85.245 192.830 85.290 ;
        RECT 195.835 85.245 195.975 85.740 ;
        RECT 196.205 85.725 196.525 85.985 ;
        RECT 196.665 85.725 196.985 85.985 ;
        RECT 201.355 85.970 201.495 86.125 ;
        RECT 201.280 85.740 201.570 85.970 ;
        RECT 201.725 85.925 202.045 85.985 ;
        RECT 202.200 85.925 202.490 85.970 ;
        RECT 201.725 85.785 202.490 85.925 ;
        RECT 203.655 85.925 203.795 86.465 ;
        RECT 210.005 86.265 210.325 86.325 ;
        RECT 205.495 86.125 210.325 86.265 ;
        RECT 205.495 85.970 205.635 86.125 ;
        RECT 210.005 86.065 210.325 86.125 ;
        RECT 210.555 85.985 210.695 86.465 ;
        RECT 212.765 86.265 213.085 86.325 ;
        RECT 211.935 86.125 213.085 86.265 ;
        RECT 204.040 85.925 204.330 85.970 ;
        RECT 203.655 85.785 204.330 85.925 ;
        RECT 201.355 85.305 201.495 85.740 ;
        RECT 201.725 85.725 202.045 85.785 ;
        RECT 202.200 85.740 202.490 85.785 ;
        RECT 204.040 85.740 204.330 85.785 ;
        RECT 204.960 85.740 205.250 85.970 ;
        RECT 205.420 85.740 205.710 85.970 ;
        RECT 203.120 85.585 203.410 85.630 ;
        RECT 205.035 85.585 205.175 85.740 ;
        RECT 205.865 85.725 206.185 85.985 ;
        RECT 208.625 85.925 208.945 85.985 ;
        RECT 209.100 85.925 209.390 85.970 ;
        RECT 208.625 85.785 209.390 85.925 ;
        RECT 208.625 85.725 208.945 85.785 ;
        RECT 209.100 85.740 209.390 85.785 ;
        RECT 210.465 85.725 210.785 85.985 ;
        RECT 211.935 85.970 212.075 86.125 ;
        RECT 212.765 86.065 213.085 86.125 ;
        RECT 223.345 86.265 223.665 86.325 ;
        RECT 226.565 86.265 226.885 86.325 ;
        RECT 242.755 86.265 242.895 86.745 ;
        RECT 244.505 86.605 244.825 86.665 ;
        RECT 247.725 86.605 248.045 86.665 ;
        RECT 244.505 86.465 248.045 86.605 ;
        RECT 244.505 86.405 244.825 86.465 ;
        RECT 247.725 86.405 248.045 86.465 ;
        RECT 248.645 86.265 248.965 86.325 ;
        RECT 223.345 86.125 242.895 86.265 ;
        RECT 244.595 86.125 248.965 86.265 ;
        RECT 249.170 86.265 249.310 86.805 ;
        RECT 250.485 86.745 250.805 87.005 ;
        RECT 258.305 86.945 258.625 87.005 ;
        RECT 276.245 86.945 276.565 87.005 ;
        RECT 258.305 86.805 276.565 86.945 ;
        RECT 258.305 86.745 258.625 86.805 ;
        RECT 276.245 86.745 276.565 86.805 ;
        RECT 286.825 86.745 287.145 87.005 ;
        RECT 297.865 86.945 298.185 87.005 ;
        RECT 308.920 86.945 309.210 86.990 ;
        RECT 297.865 86.805 309.210 86.945 ;
        RECT 297.865 86.745 298.185 86.805 ;
        RECT 308.920 86.760 309.210 86.805 ;
        RECT 252.325 86.605 252.645 86.665 ;
        RECT 267.505 86.605 267.825 86.665 ;
        RECT 252.325 86.465 267.825 86.605 ;
        RECT 252.325 86.405 252.645 86.465 ;
        RECT 267.505 86.405 267.825 86.465 ;
        RECT 295.530 86.605 295.820 86.650 ;
        RECT 297.420 86.605 297.710 86.650 ;
        RECT 300.540 86.605 300.830 86.650 ;
        RECT 295.530 86.465 300.830 86.605 ;
        RECT 295.530 86.420 295.820 86.465 ;
        RECT 297.420 86.420 297.710 86.465 ;
        RECT 300.540 86.420 300.830 86.465 ;
        RECT 306.620 86.605 306.910 86.650 ;
        RECT 310.285 86.605 310.605 86.665 ;
        RECT 306.620 86.465 310.605 86.605 ;
        RECT 306.620 86.420 306.910 86.465 ;
        RECT 310.285 86.405 310.605 86.465 ;
        RECT 256.465 86.265 256.785 86.325 ;
        RECT 260.605 86.265 260.925 86.325 ;
        RECT 249.170 86.125 260.925 86.265 ;
        RECT 223.345 86.065 223.665 86.125 ;
        RECT 226.565 86.065 226.885 86.125 ;
        RECT 211.400 85.740 211.690 85.970 ;
        RECT 211.860 85.740 212.150 85.970 ;
        RECT 208.180 85.585 208.470 85.630 ;
        RECT 203.120 85.445 205.175 85.585 ;
        RECT 205.495 85.445 208.470 85.585 ;
        RECT 203.120 85.400 203.410 85.445 ;
        RECT 192.540 85.105 195.975 85.245 ;
        RECT 198.060 85.245 198.350 85.290 ;
        RECT 198.505 85.245 198.825 85.305 ;
        RECT 198.060 85.105 198.825 85.245 ;
        RECT 192.540 85.060 192.830 85.105 ;
        RECT 198.060 85.060 198.350 85.105 ;
        RECT 198.505 85.045 198.825 85.105 ;
        RECT 201.265 85.245 201.585 85.305 ;
        RECT 205.495 85.245 205.635 85.445 ;
        RECT 208.180 85.400 208.470 85.445 ;
        RECT 210.020 85.585 210.310 85.630 ;
        RECT 211.475 85.585 211.615 85.740 ;
        RECT 212.305 85.725 212.625 85.985 ;
        RECT 220.125 85.925 220.445 85.985 ;
        RECT 228.865 85.925 229.185 85.985 ;
        RECT 220.125 85.785 229.185 85.925 ;
        RECT 220.125 85.725 220.445 85.785 ;
        RECT 228.865 85.725 229.185 85.785 ;
        RECT 233.005 85.925 233.325 85.985 ;
        RECT 244.595 85.970 244.735 86.125 ;
        RECT 248.645 86.065 248.965 86.125 ;
        RECT 256.465 86.065 256.785 86.125 ;
        RECT 260.605 86.065 260.925 86.125 ;
        RECT 269.360 86.265 269.650 86.310 ;
        RECT 269.805 86.265 270.125 86.325 ;
        RECT 269.360 86.125 270.125 86.265 ;
        RECT 269.360 86.080 269.650 86.125 ;
        RECT 269.805 86.065 270.125 86.125 ;
        RECT 283.605 86.265 283.925 86.325 ;
        RECT 306.145 86.265 306.465 86.325 ;
        RECT 283.605 86.125 289.355 86.265 ;
        RECT 283.605 86.065 283.925 86.125 ;
        RECT 244.520 85.925 244.810 85.970 ;
        RECT 233.005 85.785 244.810 85.925 ;
        RECT 233.005 85.725 233.325 85.785 ;
        RECT 244.520 85.740 244.810 85.785 ;
        RECT 245.900 85.925 246.190 85.970 ;
        RECT 247.280 85.925 247.570 85.970 ;
        RECT 247.725 85.925 248.045 85.985 ;
        RECT 245.900 85.785 248.045 85.925 ;
        RECT 245.900 85.740 246.190 85.785 ;
        RECT 247.280 85.740 247.570 85.785 ;
        RECT 247.725 85.725 248.045 85.785 ;
        RECT 249.105 85.725 249.425 85.985 ;
        RECT 249.705 85.925 249.995 85.970 ;
        RECT 273.040 85.925 273.330 85.970 ;
        RECT 286.380 85.925 286.670 85.970 ;
        RECT 287.285 85.925 287.605 85.985 ;
        RECT 249.705 85.785 269.805 85.925 ;
        RECT 249.705 85.740 249.995 85.785 ;
        RECT 210.020 85.445 211.615 85.585 ;
        RECT 213.225 85.585 213.545 85.645 ;
        RECT 225.185 85.585 225.505 85.645 ;
        RECT 241.285 85.585 241.605 85.645 ;
        RECT 253.245 85.585 253.565 85.645 ;
        RECT 213.225 85.445 228.635 85.585 ;
        RECT 210.020 85.400 210.310 85.445 ;
        RECT 213.225 85.385 213.545 85.445 ;
        RECT 225.185 85.385 225.505 85.445 ;
        RECT 228.495 85.305 228.635 85.445 ;
        RECT 241.285 85.445 253.565 85.585 ;
        RECT 241.285 85.385 241.605 85.445 ;
        RECT 253.245 85.385 253.565 85.445 ;
        RECT 255.085 85.585 255.405 85.645 ;
        RECT 266.585 85.585 266.905 85.645 ;
        RECT 255.085 85.445 266.905 85.585 ;
        RECT 269.665 85.585 269.805 85.785 ;
        RECT 273.040 85.785 287.605 85.925 ;
        RECT 273.040 85.740 273.330 85.785 ;
        RECT 286.380 85.740 286.670 85.785 ;
        RECT 287.285 85.725 287.605 85.785 ;
        RECT 287.745 85.725 288.065 85.985 ;
        RECT 289.215 85.970 289.355 86.125 ;
        RECT 306.145 86.125 308.215 86.265 ;
        RECT 306.145 86.065 306.465 86.125 ;
        RECT 289.140 85.740 289.430 85.970 ;
        RECT 294.645 85.725 294.965 85.985 ;
        RECT 295.125 85.925 295.415 85.970 ;
        RECT 296.960 85.925 297.250 85.970 ;
        RECT 300.540 85.925 300.830 85.970 ;
        RECT 295.125 85.785 300.830 85.925 ;
        RECT 295.125 85.740 295.415 85.785 ;
        RECT 296.960 85.740 297.250 85.785 ;
        RECT 300.540 85.740 300.830 85.785 ;
        RECT 282.700 85.585 282.990 85.630 ;
        RECT 283.605 85.585 283.925 85.645 ;
        RECT 294.735 85.585 294.875 85.725 ;
        RECT 269.665 85.445 282.455 85.585 ;
        RECT 255.085 85.385 255.405 85.445 ;
        RECT 266.585 85.385 266.905 85.445 ;
        RECT 201.265 85.105 205.635 85.245 ;
        RECT 207.260 85.245 207.550 85.290 ;
        RECT 207.705 85.245 208.025 85.305 ;
        RECT 207.260 85.105 208.025 85.245 ;
        RECT 201.265 85.045 201.585 85.105 ;
        RECT 207.260 85.060 207.550 85.105 ;
        RECT 207.705 85.045 208.025 85.105 ;
        RECT 213.700 85.245 213.990 85.290 ;
        RECT 216.445 85.245 216.765 85.305 ;
        RECT 213.700 85.105 216.765 85.245 ;
        RECT 213.700 85.060 213.990 85.105 ;
        RECT 216.445 85.045 216.765 85.105 ;
        RECT 228.405 85.045 228.725 85.305 ;
        RECT 244.965 85.245 245.285 85.305 ;
        RECT 250.025 85.245 250.345 85.305 ;
        RECT 270.265 85.245 270.585 85.305 ;
        RECT 244.965 85.105 270.585 85.245 ;
        RECT 282.315 85.245 282.455 85.445 ;
        RECT 282.700 85.445 294.875 85.585 ;
        RECT 295.565 85.585 295.885 85.645 ;
        RECT 296.040 85.585 296.330 85.630 ;
        RECT 295.565 85.445 296.330 85.585 ;
        RECT 282.700 85.400 282.990 85.445 ;
        RECT 283.605 85.385 283.925 85.445 ;
        RECT 295.565 85.385 295.885 85.445 ;
        RECT 296.040 85.400 296.330 85.445 ;
        RECT 298.320 85.585 298.970 85.630 ;
        RECT 299.705 85.585 300.025 85.645 ;
        RECT 301.620 85.630 301.910 85.945 ;
        RECT 307.525 85.725 307.845 85.985 ;
        RECT 308.075 85.970 308.215 86.125 ;
        RECT 308.000 85.740 308.290 85.970 ;
        RECT 301.620 85.585 302.210 85.630 ;
        RECT 298.320 85.445 302.210 85.585 ;
        RECT 298.320 85.400 298.970 85.445 ;
        RECT 299.705 85.385 300.025 85.445 ;
        RECT 301.920 85.400 302.210 85.445 ;
        RECT 288.680 85.245 288.970 85.290 ;
        RECT 302.925 85.245 303.245 85.305 ;
        RECT 303.400 85.245 303.690 85.290 ;
        RECT 282.315 85.105 303.690 85.245 ;
        RECT 244.965 85.045 245.285 85.105 ;
        RECT 250.025 85.045 250.345 85.105 ;
        RECT 270.265 85.045 270.585 85.105 ;
        RECT 288.680 85.060 288.970 85.105 ;
        RECT 302.925 85.045 303.245 85.105 ;
        RECT 303.400 85.060 303.690 85.105 ;
        RECT 162.095 84.425 311.135 84.905 ;
        RECT 166.305 84.225 166.625 84.285 ;
        RECT 172.745 84.225 173.065 84.285 ;
        RECT 175.520 84.225 175.810 84.270 ;
        RECT 212.305 84.225 212.625 84.285 ;
        RECT 230.245 84.225 230.565 84.285 ;
        RECT 251.420 84.225 251.710 84.270 ;
        RECT 166.305 84.085 216.215 84.225 ;
        RECT 166.305 84.025 166.625 84.085 ;
        RECT 172.745 84.025 173.065 84.085 ;
        RECT 175.520 84.040 175.810 84.085 ;
        RECT 212.305 84.025 212.625 84.085 ;
        RECT 167.685 83.885 168.005 83.945 ;
        RECT 166.855 83.745 168.005 83.885 ;
        RECT 166.855 83.590 166.995 83.745 ;
        RECT 167.685 83.685 168.005 83.745 ;
        RECT 170.440 83.885 171.090 83.930 ;
        RECT 174.040 83.885 174.330 83.930 ;
        RECT 176.885 83.885 177.205 83.945 ;
        RECT 170.440 83.745 177.205 83.885 ;
        RECT 170.440 83.700 171.090 83.745 ;
        RECT 173.740 83.700 174.330 83.745 ;
        RECT 166.780 83.360 167.070 83.590 ;
        RECT 167.245 83.545 167.535 83.590 ;
        RECT 169.080 83.545 169.370 83.590 ;
        RECT 172.660 83.545 172.950 83.590 ;
        RECT 167.245 83.405 172.950 83.545 ;
        RECT 167.245 83.360 167.535 83.405 ;
        RECT 169.080 83.360 169.370 83.405 ;
        RECT 172.660 83.360 172.950 83.405 ;
        RECT 173.740 83.385 174.030 83.700 ;
        RECT 176.885 83.685 177.205 83.745 ;
        RECT 184.720 83.885 185.010 83.930 ;
        RECT 186.085 83.885 186.405 83.945 ;
        RECT 184.720 83.745 186.405 83.885 ;
        RECT 184.720 83.700 185.010 83.745 ;
        RECT 186.085 83.685 186.405 83.745 ;
        RECT 188.845 83.685 189.165 83.945 ;
        RECT 193.445 83.885 193.765 83.945 ;
        RECT 200.360 83.885 200.650 83.930 ;
        RECT 208.640 83.885 208.930 83.930 ;
        RECT 193.445 83.745 208.930 83.885 ;
        RECT 193.445 83.685 193.765 83.745 ;
        RECT 200.360 83.700 200.650 83.745 ;
        RECT 208.640 83.700 208.930 83.745 ;
        RECT 210.465 83.885 210.785 83.945 ;
        RECT 210.465 83.745 214.375 83.885 ;
        RECT 210.465 83.685 210.785 83.745 ;
        RECT 185.640 83.545 185.930 83.590 ;
        RECT 189.765 83.545 190.085 83.605 ;
        RECT 185.640 83.405 190.085 83.545 ;
        RECT 185.640 83.360 185.930 83.405 ;
        RECT 189.765 83.345 190.085 83.405 ;
        RECT 192.985 83.545 193.305 83.605 ;
        RECT 196.220 83.545 196.510 83.590 ;
        RECT 192.985 83.405 196.510 83.545 ;
        RECT 192.985 83.345 193.305 83.405 ;
        RECT 196.220 83.360 196.510 83.405 ;
        RECT 205.880 83.545 206.170 83.590 ;
        RECT 211.845 83.545 212.165 83.605 ;
        RECT 214.235 83.590 214.375 83.745 ;
        RECT 212.320 83.545 212.610 83.590 ;
        RECT 205.880 83.405 212.610 83.545 ;
        RECT 205.880 83.360 206.170 83.405 ;
        RECT 211.845 83.345 212.165 83.405 ;
        RECT 212.320 83.360 212.610 83.405 ;
        RECT 214.160 83.360 214.450 83.590 ;
        RECT 215.065 83.345 215.385 83.605 ;
        RECT 216.075 83.590 216.215 84.085 ;
        RECT 227.115 84.085 230.565 84.225 ;
        RECT 227.115 83.590 227.255 84.085 ;
        RECT 230.245 84.025 230.565 84.085 ;
        RECT 240.915 84.085 251.710 84.225 ;
        RECT 227.485 83.885 227.805 83.945 ;
        RECT 240.915 83.930 241.055 84.085 ;
        RECT 251.420 84.040 251.710 84.085 ;
        RECT 302.005 84.225 302.325 84.285 ;
        RECT 304.780 84.225 305.070 84.270 ;
        RECT 302.005 84.085 305.070 84.225 ;
        RECT 302.005 84.025 302.325 84.085 ;
        RECT 304.780 84.040 305.070 84.085 ;
        RECT 240.840 83.885 241.130 83.930 ;
        RECT 227.485 83.745 241.130 83.885 ;
        RECT 227.485 83.685 227.805 83.745 ;
        RECT 240.840 83.700 241.130 83.745 ;
        RECT 242.665 83.885 242.985 83.945 ;
        RECT 244.060 83.885 244.350 83.930 ;
        RECT 242.665 83.745 244.350 83.885 ;
        RECT 242.665 83.685 242.985 83.745 ;
        RECT 244.060 83.700 244.350 83.745 ;
        RECT 244.505 83.685 244.825 83.945 ;
        RECT 248.185 83.885 248.505 83.945 ;
        RECT 252.340 83.885 252.630 83.930 ;
        RECT 246.435 83.745 252.630 83.885 ;
        RECT 246.435 83.605 246.575 83.745 ;
        RECT 248.185 83.685 248.505 83.745 ;
        RECT 252.340 83.700 252.630 83.745 ;
        RECT 253.245 83.885 253.565 83.945 ;
        RECT 257.385 83.885 257.705 83.945 ;
        RECT 253.245 83.745 257.705 83.885 ;
        RECT 253.245 83.685 253.565 83.745 ;
        RECT 257.385 83.685 257.705 83.745 ;
        RECT 276.245 83.885 276.565 83.945 ;
        RECT 279.020 83.885 279.310 83.930 ;
        RECT 276.245 83.745 279.310 83.885 ;
        RECT 276.245 83.685 276.565 83.745 ;
        RECT 279.020 83.700 279.310 83.745 ;
        RECT 296.945 83.885 297.265 83.945 ;
        RECT 299.705 83.930 300.025 83.945 ;
        RECT 297.420 83.885 297.710 83.930 ;
        RECT 296.945 83.745 297.710 83.885 ;
        RECT 296.945 83.685 297.265 83.745 ;
        RECT 297.420 83.700 297.710 83.745 ;
        RECT 299.700 83.885 300.350 83.930 ;
        RECT 303.300 83.885 303.590 83.930 ;
        RECT 299.700 83.745 303.590 83.885 ;
        RECT 299.700 83.700 300.350 83.745 ;
        RECT 303.000 83.700 303.590 83.745 ;
        RECT 299.705 83.685 300.025 83.700 ;
        RECT 215.540 83.360 215.830 83.590 ;
        RECT 216.000 83.360 216.290 83.590 ;
        RECT 227.040 83.360 227.330 83.590 ;
        RECT 168.160 83.205 168.450 83.250 ;
        RECT 170.905 83.205 171.225 83.265 ;
        RECT 168.160 83.065 171.225 83.205 ;
        RECT 168.160 83.020 168.450 83.065 ;
        RECT 170.905 83.005 171.225 83.065 ;
        RECT 183.785 83.205 184.105 83.265 ;
        RECT 186.560 83.205 186.850 83.250 ;
        RECT 183.785 83.065 186.850 83.205 ;
        RECT 183.785 83.005 184.105 83.065 ;
        RECT 186.560 83.020 186.850 83.065 ;
        RECT 190.685 83.005 191.005 83.265 ;
        RECT 199.885 83.205 200.205 83.265 ;
        RECT 215.615 83.205 215.755 83.360 ;
        RECT 227.945 83.345 228.265 83.605 ;
        RECT 228.405 83.345 228.725 83.605 ;
        RECT 228.880 83.360 229.170 83.590 ;
        RECT 229.325 83.545 229.645 83.605 ;
        RECT 243.585 83.590 243.905 83.605 ;
        RECT 242.220 83.545 242.510 83.590 ;
        RECT 243.575 83.545 243.905 83.590 ;
        RECT 229.325 83.405 242.510 83.545 ;
        RECT 243.390 83.405 243.905 83.545 ;
        RECT 199.885 83.065 215.755 83.205 ;
        RECT 199.885 83.005 200.205 83.065 ;
        RECT 217.365 83.005 217.685 83.265 ;
        RECT 167.650 82.865 167.940 82.910 ;
        RECT 169.540 82.865 169.830 82.910 ;
        RECT 172.660 82.865 172.950 82.910 ;
        RECT 167.650 82.725 172.950 82.865 ;
        RECT 167.650 82.680 167.940 82.725 ;
        RECT 169.540 82.680 169.830 82.725 ;
        RECT 172.660 82.680 172.950 82.725 ;
        RECT 206.785 82.865 207.105 82.925 ;
        RECT 226.565 82.865 226.885 82.925 ;
        RECT 228.950 82.865 229.090 83.360 ;
        RECT 229.325 83.345 229.645 83.405 ;
        RECT 242.220 83.360 242.510 83.405 ;
        RECT 243.575 83.360 243.905 83.405 ;
        RECT 242.295 83.205 242.435 83.360 ;
        RECT 243.585 83.345 243.905 83.360 ;
        RECT 244.965 83.590 245.285 83.605 ;
        RECT 244.965 83.360 245.450 83.590 ;
        RECT 245.900 83.545 246.190 83.590 ;
        RECT 246.345 83.545 246.665 83.605 ;
        RECT 245.900 83.405 246.665 83.545 ;
        RECT 245.900 83.360 246.190 83.405 ;
        RECT 244.965 83.345 245.285 83.360 ;
        RECT 246.345 83.345 246.665 83.405 ;
        RECT 247.265 83.345 247.585 83.605 ;
        RECT 248.645 83.345 248.965 83.605 ;
        RECT 250.485 83.345 250.805 83.605 ;
        RECT 256.925 83.545 257.245 83.605 ;
        RECT 260.620 83.545 260.910 83.590 ;
        RECT 256.925 83.405 260.910 83.545 ;
        RECT 256.925 83.345 257.245 83.405 ;
        RECT 260.620 83.360 260.910 83.405 ;
        RECT 261.065 83.545 261.385 83.605 ;
        RECT 261.540 83.545 261.830 83.590 ;
        RECT 261.065 83.405 261.830 83.545 ;
        RECT 261.065 83.345 261.385 83.405 ;
        RECT 261.540 83.360 261.830 83.405 ;
        RECT 262.000 83.545 262.290 83.590 ;
        RECT 265.205 83.545 265.525 83.605 ;
        RECT 262.000 83.405 265.525 83.545 ;
        RECT 262.000 83.360 262.290 83.405 ;
        RECT 265.205 83.345 265.525 83.405 ;
        RECT 266.585 83.345 266.905 83.605 ;
        RECT 269.805 83.345 270.125 83.605 ;
        RECT 278.085 83.345 278.405 83.605 ;
        RECT 283.605 83.345 283.925 83.605 ;
        RECT 293.740 83.545 294.030 83.590 ;
        RECT 295.105 83.545 295.425 83.605 ;
        RECT 293.740 83.405 295.425 83.545 ;
        RECT 293.740 83.360 294.030 83.405 ;
        RECT 295.105 83.345 295.425 83.405 ;
        RECT 296.025 83.345 296.345 83.605 ;
        RECT 296.505 83.545 296.795 83.590 ;
        RECT 298.340 83.545 298.630 83.590 ;
        RECT 301.920 83.545 302.210 83.590 ;
        RECT 296.505 83.405 302.210 83.545 ;
        RECT 296.505 83.360 296.795 83.405 ;
        RECT 298.340 83.360 298.630 83.405 ;
        RECT 301.920 83.360 302.210 83.405 ;
        RECT 303.000 83.385 303.290 83.700 ;
        RECT 247.725 83.205 248.045 83.265 ;
        RECT 242.295 83.065 248.045 83.205 ;
        RECT 247.725 83.005 248.045 83.065 ;
        RECT 248.185 83.005 248.505 83.265 ;
        RECT 263.365 83.205 263.685 83.265 ;
        RECT 265.680 83.205 265.970 83.250 ;
        RECT 263.365 83.065 265.970 83.205 ;
        RECT 263.365 83.005 263.685 83.065 ;
        RECT 265.680 83.020 265.970 83.065 ;
        RECT 274.405 83.205 274.725 83.265 ;
        RECT 277.180 83.205 277.470 83.250 ;
        RECT 274.405 83.065 277.470 83.205 ;
        RECT 274.405 83.005 274.725 83.065 ;
        RECT 277.180 83.020 277.470 83.065 ;
        RECT 206.785 82.725 226.335 82.865 ;
        RECT 206.785 82.665 207.105 82.725 ;
        RECT 226.195 82.525 226.335 82.725 ;
        RECT 226.565 82.725 229.090 82.865 ;
        RECT 229.325 82.865 229.645 82.925 ;
        RECT 241.760 82.865 242.050 82.910 ;
        RECT 259.685 82.865 260.005 82.925 ;
        RECT 261.985 82.865 262.305 82.925 ;
        RECT 229.325 82.725 247.955 82.865 ;
        RECT 226.565 82.665 226.885 82.725 ;
        RECT 229.325 82.665 229.645 82.725 ;
        RECT 241.760 82.680 242.050 82.725 ;
        RECT 227.945 82.525 228.265 82.585 ;
        RECT 226.195 82.385 228.265 82.525 ;
        RECT 227.945 82.325 228.265 82.385 ;
        RECT 229.800 82.525 230.090 82.570 ;
        RECT 233.465 82.525 233.785 82.585 ;
        RECT 229.800 82.385 233.785 82.525 ;
        RECT 229.800 82.340 230.090 82.385 ;
        RECT 233.465 82.325 233.785 82.385 ;
        RECT 241.285 82.325 241.605 82.585 ;
        RECT 242.205 82.525 242.525 82.585 ;
        RECT 242.680 82.525 242.970 82.570 ;
        RECT 242.205 82.385 242.970 82.525 ;
        RECT 242.205 82.325 242.525 82.385 ;
        RECT 242.680 82.340 242.970 82.385 ;
        RECT 246.360 82.525 246.650 82.570 ;
        RECT 247.265 82.525 247.585 82.585 ;
        RECT 246.360 82.385 247.585 82.525 ;
        RECT 247.815 82.525 247.955 82.725 ;
        RECT 259.685 82.725 262.305 82.865 ;
        RECT 259.685 82.665 260.005 82.725 ;
        RECT 261.985 82.665 262.305 82.725 ;
        RECT 296.910 82.865 297.200 82.910 ;
        RECT 298.800 82.865 299.090 82.910 ;
        RECT 301.920 82.865 302.210 82.910 ;
        RECT 296.910 82.725 302.210 82.865 ;
        RECT 296.910 82.680 297.200 82.725 ;
        RECT 298.800 82.680 299.090 82.725 ;
        RECT 301.920 82.680 302.210 82.725 ;
        RECT 249.565 82.525 249.885 82.585 ;
        RECT 247.815 82.385 249.885 82.525 ;
        RECT 246.360 82.340 246.650 82.385 ;
        RECT 247.265 82.325 247.585 82.385 ;
        RECT 249.565 82.325 249.885 82.385 ;
        RECT 260.605 82.325 260.925 82.585 ;
        RECT 262.905 82.325 263.225 82.585 ;
        RECT 267.520 82.525 267.810 82.570 ;
        RECT 269.345 82.525 269.665 82.585 ;
        RECT 267.520 82.385 269.665 82.525 ;
        RECT 267.520 82.340 267.810 82.385 ;
        RECT 269.345 82.325 269.665 82.385 ;
        RECT 162.095 81.705 311.135 82.185 ;
        RECT 170.905 81.305 171.225 81.565 ;
        RECT 204.945 81.505 205.265 81.565 ;
        RECT 212.765 81.505 213.085 81.565 ;
        RECT 204.945 81.365 213.085 81.505 ;
        RECT 204.945 81.305 205.265 81.365 ;
        RECT 212.765 81.305 213.085 81.365 ;
        RECT 218.300 81.505 218.590 81.550 ;
        RECT 223.345 81.505 223.665 81.565 ;
        RECT 218.300 81.365 223.665 81.505 ;
        RECT 218.300 81.320 218.590 81.365 ;
        RECT 223.345 81.305 223.665 81.365 ;
        RECT 224.740 81.505 225.030 81.550 ;
        RECT 233.005 81.505 233.325 81.565 ;
        RECT 242.205 81.505 242.525 81.565 ;
        RECT 224.740 81.365 233.325 81.505 ;
        RECT 224.740 81.320 225.030 81.365 ;
        RECT 233.005 81.305 233.325 81.365 ;
        RECT 234.475 81.365 242.525 81.505 ;
        RECT 174.125 81.165 174.445 81.225 ;
        RECT 175.520 81.165 175.810 81.210 ;
        RECT 187.005 81.165 187.325 81.225 ;
        RECT 194.365 81.165 194.685 81.225 ;
        RECT 174.125 81.025 175.810 81.165 ;
        RECT 174.125 80.965 174.445 81.025 ;
        RECT 175.520 80.980 175.810 81.025 ;
        RECT 178.355 81.025 194.685 81.165 ;
        RECT 172.285 80.825 172.605 80.885 ;
        RECT 173.680 80.825 173.970 80.870 ;
        RECT 172.285 80.685 173.970 80.825 ;
        RECT 172.285 80.625 172.605 80.685 ;
        RECT 173.680 80.640 173.970 80.685 ;
        RECT 175.045 80.825 175.365 80.885 ;
        RECT 178.355 80.825 178.495 81.025 ;
        RECT 187.005 80.965 187.325 81.025 ;
        RECT 194.365 80.965 194.685 81.025 ;
        RECT 194.840 81.165 195.130 81.210 ;
        RECT 195.745 81.165 196.065 81.225 ;
        RECT 229.325 81.165 229.645 81.225 ;
        RECT 233.925 81.165 234.245 81.225 ;
        RECT 194.840 81.025 196.065 81.165 ;
        RECT 194.840 80.980 195.130 81.025 ;
        RECT 195.745 80.965 196.065 81.025 ;
        RECT 213.315 81.025 229.645 81.165 ;
        RECT 175.045 80.685 178.495 80.825 ;
        RECT 178.740 80.825 179.030 80.870 ;
        RECT 179.645 80.825 179.965 80.885 ;
        RECT 178.740 80.685 179.965 80.825 ;
        RECT 175.045 80.625 175.365 80.685 ;
        RECT 178.740 80.640 179.030 80.685 ;
        RECT 179.645 80.625 179.965 80.685 ;
        RECT 184.245 80.825 184.565 80.885 ;
        RECT 194.455 80.825 194.595 80.965 ;
        RECT 196.680 80.825 196.970 80.870 ;
        RECT 207.245 80.825 207.565 80.885 ;
        RECT 213.315 80.825 213.455 81.025 ;
        RECT 229.325 80.965 229.645 81.025 ;
        RECT 230.795 81.025 234.245 81.165 ;
        RECT 223.805 80.825 224.125 80.885 ;
        RECT 226.105 80.825 226.425 80.885 ;
        RECT 184.245 80.685 192.295 80.825 ;
        RECT 194.455 80.685 196.435 80.825 ;
        RECT 184.245 80.625 184.565 80.685 ;
        RECT 173.220 80.485 173.510 80.530 ;
        RECT 185.165 80.485 185.485 80.545 ;
        RECT 173.220 80.345 185.485 80.485 ;
        RECT 173.220 80.300 173.510 80.345 ;
        RECT 185.165 80.285 185.485 80.345 ;
        RECT 191.605 80.285 191.925 80.545 ;
        RECT 192.155 80.485 192.295 80.685 ;
        RECT 194.380 80.485 194.670 80.530 ;
        RECT 192.155 80.345 194.670 80.485 ;
        RECT 194.380 80.300 194.670 80.345 ;
        RECT 195.285 80.485 195.605 80.545 ;
        RECT 195.760 80.485 196.050 80.530 ;
        RECT 195.285 80.345 196.050 80.485 ;
        RECT 196.295 80.485 196.435 80.685 ;
        RECT 196.680 80.685 207.565 80.825 ;
        RECT 196.680 80.640 196.970 80.685 ;
        RECT 207.245 80.625 207.565 80.685 ;
        RECT 208.255 80.685 209.315 80.825 ;
        RECT 204.945 80.485 205.265 80.545 ;
        RECT 196.295 80.345 205.265 80.485 ;
        RECT 195.285 80.285 195.605 80.345 ;
        RECT 195.760 80.300 196.050 80.345 ;
        RECT 204.945 80.285 205.265 80.345 ;
        RECT 205.880 80.485 206.170 80.530 ;
        RECT 208.255 80.485 208.395 80.685 ;
        RECT 205.880 80.345 208.395 80.485 ;
        RECT 205.880 80.300 206.170 80.345 ;
        RECT 172.745 79.945 173.065 80.205 ;
        RECT 176.425 80.145 176.745 80.205 ;
        RECT 177.820 80.145 178.110 80.190 ;
        RECT 180.105 80.145 180.425 80.205 ;
        RECT 176.425 80.005 180.425 80.145 ;
        RECT 176.425 79.945 176.745 80.005 ;
        RECT 177.820 79.960 178.110 80.005 ;
        RECT 180.105 79.945 180.425 80.005 ;
        RECT 182.865 80.145 183.185 80.205 ;
        RECT 193.905 80.145 194.225 80.205 ;
        RECT 205.955 80.145 206.095 80.300 ;
        RECT 208.625 80.285 208.945 80.545 ;
        RECT 209.175 80.485 209.315 80.685 ;
        RECT 212.395 80.685 213.455 80.825 ;
        RECT 213.775 80.685 224.125 80.825 ;
        RECT 211.860 80.485 212.150 80.530 ;
        RECT 212.395 80.485 212.535 80.685 ;
        RECT 209.175 80.345 212.535 80.485 ;
        RECT 212.765 80.485 213.085 80.545 ;
        RECT 213.775 80.485 213.915 80.685 ;
        RECT 223.805 80.625 224.125 80.685 ;
        RECT 224.355 80.685 229.990 80.825 ;
        RECT 212.765 80.345 213.915 80.485 ;
        RECT 211.860 80.300 212.150 80.345 ;
        RECT 212.765 80.285 213.085 80.345 ;
        RECT 215.065 80.285 215.385 80.545 ;
        RECT 224.355 80.485 224.495 80.685 ;
        RECT 226.105 80.625 226.425 80.685 ;
        RECT 229.850 80.530 229.990 80.685 ;
        RECT 215.615 80.345 224.495 80.485 ;
        RECT 206.325 80.145 206.645 80.205 ;
        RECT 182.865 80.005 190.915 80.145 ;
        RECT 182.865 79.945 183.185 80.005 ;
        RECT 175.965 79.805 176.285 79.865 ;
        RECT 177.360 79.805 177.650 79.850 ;
        RECT 175.965 79.665 177.650 79.805 ;
        RECT 190.775 79.805 190.915 80.005 ;
        RECT 193.905 80.005 206.645 80.145 ;
        RECT 193.905 79.945 194.225 80.005 ;
        RECT 206.325 79.945 206.645 80.005 ;
        RECT 208.165 80.145 208.485 80.205 ;
        RECT 211.400 80.145 211.690 80.190 ;
        RECT 215.615 80.145 215.755 80.345 ;
        RECT 229.775 80.300 230.065 80.530 ;
        RECT 208.165 80.005 215.755 80.145 ;
        RECT 223.805 80.145 224.125 80.205 ;
        RECT 227.485 80.145 227.805 80.205 ;
        RECT 223.805 80.005 227.805 80.145 ;
        RECT 208.165 79.945 208.485 80.005 ;
        RECT 211.400 79.960 211.690 80.005 ;
        RECT 223.805 79.945 224.125 80.005 ;
        RECT 227.485 79.945 227.805 80.005 ;
        RECT 197.585 79.805 197.905 79.865 ;
        RECT 220.585 79.805 220.905 79.865 ;
        RECT 190.775 79.665 220.905 79.805 ;
        RECT 175.965 79.605 176.285 79.665 ;
        RECT 177.360 79.620 177.650 79.665 ;
        RECT 197.585 79.605 197.905 79.665 ;
        RECT 220.585 79.605 220.905 79.665 ;
        RECT 224.725 79.605 225.045 79.865 ;
        RECT 225.660 79.805 225.950 79.850 ;
        RECT 226.565 79.805 226.885 79.865 ;
        RECT 225.660 79.665 226.885 79.805 ;
        RECT 225.660 79.620 225.950 79.665 ;
        RECT 226.565 79.605 226.885 79.665 ;
        RECT 228.405 79.805 228.725 79.865 ;
        RECT 228.880 79.805 229.170 79.850 ;
        RECT 228.405 79.665 229.170 79.805 ;
        RECT 229.850 79.805 229.990 80.300 ;
        RECT 230.245 80.285 230.565 80.545 ;
        RECT 230.795 80.530 230.935 81.025 ;
        RECT 233.925 80.965 234.245 81.025 ;
        RECT 234.475 80.825 234.615 81.365 ;
        RECT 242.205 81.305 242.525 81.365 ;
        RECT 243.585 81.505 243.905 81.565 ;
        RECT 246.805 81.505 247.125 81.565 ;
        RECT 243.585 81.365 247.125 81.505 ;
        RECT 243.585 81.305 243.905 81.365 ;
        RECT 246.805 81.305 247.125 81.365 ;
        RECT 247.725 81.305 248.045 81.565 ;
        RECT 248.645 81.505 248.965 81.565 ;
        RECT 248.645 81.365 256.005 81.505 ;
        RECT 248.645 81.305 248.965 81.365 ;
        RECT 240.365 81.165 240.685 81.225 ;
        RECT 255.085 81.165 255.405 81.225 ;
        RECT 240.365 81.025 255.405 81.165 ;
        RECT 255.865 81.165 256.005 81.365 ;
        RECT 256.925 81.305 257.245 81.565 ;
        RECT 264.760 81.505 265.050 81.550 ;
        RECT 267.980 81.505 268.270 81.550 ;
        RECT 264.760 81.365 268.270 81.505 ;
        RECT 264.760 81.320 265.050 81.365 ;
        RECT 267.980 81.320 268.270 81.365 ;
        RECT 270.265 81.505 270.585 81.565 ;
        RECT 283.605 81.505 283.925 81.565 ;
        RECT 270.265 81.365 283.925 81.505 ;
        RECT 270.265 81.305 270.585 81.365 ;
        RECT 283.605 81.305 283.925 81.365 ;
        RECT 286.365 81.505 286.685 81.565 ;
        RECT 306.605 81.505 306.925 81.565 ;
        RECT 286.365 81.365 306.925 81.505 ;
        RECT 286.365 81.305 286.685 81.365 ;
        RECT 306.605 81.305 306.925 81.365 ;
        RECT 257.385 81.165 257.705 81.225 ;
        RECT 255.865 81.025 257.155 81.165 ;
        RECT 240.365 80.965 240.685 81.025 ;
        RECT 255.085 80.965 255.405 81.025 ;
        RECT 246.345 80.825 246.665 80.885 ;
        RECT 256.465 80.825 256.785 80.885 ;
        RECT 232.175 80.685 234.615 80.825 ;
        RECT 242.755 80.685 246.665 80.825 ;
        RECT 230.720 80.300 231.010 80.530 ;
        RECT 231.625 80.285 231.945 80.545 ;
        RECT 232.175 80.530 232.315 80.685 ;
        RECT 232.100 80.300 232.390 80.530 ;
        RECT 233.465 80.285 233.785 80.545 ;
        RECT 234.385 80.285 234.705 80.545 ;
        RECT 234.860 80.485 235.150 80.530 ;
        RECT 235.305 80.485 235.625 80.545 ;
        RECT 234.860 80.345 235.625 80.485 ;
        RECT 234.860 80.300 235.150 80.345 ;
        RECT 235.305 80.285 235.625 80.345 ;
        RECT 239.445 80.285 239.765 80.545 ;
        RECT 240.365 80.285 240.685 80.545 ;
        RECT 240.825 80.285 241.145 80.545 ;
        RECT 241.300 80.485 241.590 80.530 ;
        RECT 241.745 80.485 242.065 80.545 ;
        RECT 242.755 80.530 242.895 80.685 ;
        RECT 246.345 80.625 246.665 80.685 ;
        RECT 247.360 80.685 256.785 80.825 ;
        RECT 243.585 80.530 243.905 80.545 ;
        RECT 241.300 80.345 242.065 80.485 ;
        RECT 241.300 80.300 241.590 80.345 ;
        RECT 241.745 80.285 242.065 80.345 ;
        RECT 242.680 80.300 242.970 80.530 ;
        RECT 243.420 80.300 243.905 80.530 ;
        RECT 243.585 80.285 243.905 80.300 ;
        RECT 244.045 80.285 244.365 80.545 ;
        RECT 245.210 80.485 245.500 80.530 ;
        RECT 247.360 80.485 247.500 80.685 ;
        RECT 256.465 80.625 256.785 80.685 ;
        RECT 257.015 80.545 257.155 81.025 ;
        RECT 257.385 81.025 260.790 81.165 ;
        RECT 257.385 80.965 257.705 81.025 ;
        RECT 245.210 80.345 247.500 80.485 ;
        RECT 245.210 80.300 245.500 80.345 ;
        RECT 249.565 80.285 249.885 80.545 ;
        RECT 252.785 80.485 253.105 80.545 ;
        RECT 254.165 80.485 254.485 80.545 ;
        RECT 252.785 80.345 254.485 80.485 ;
        RECT 252.785 80.285 253.105 80.345 ;
        RECT 254.165 80.285 254.485 80.345 ;
        RECT 255.085 80.285 255.405 80.545 ;
        RECT 255.545 80.285 255.865 80.545 ;
        RECT 256.020 80.485 256.310 80.530 ;
        RECT 256.925 80.485 257.245 80.545 ;
        RECT 257.475 80.530 257.615 80.965 ;
        RECT 260.145 80.825 260.465 80.885 ;
        RECT 258.855 80.685 260.465 80.825 ;
        RECT 260.650 80.825 260.790 81.025 ;
        RECT 261.065 80.965 261.385 81.225 ;
        RECT 266.125 80.965 266.445 81.225 ;
        RECT 279.925 81.165 280.245 81.225 ;
        RECT 280.860 81.165 281.150 81.210 ;
        RECT 292.345 81.165 292.665 81.225 ;
        RECT 294.645 81.165 294.965 81.225 ;
        RECT 279.925 81.025 281.150 81.165 ;
        RECT 279.925 80.965 280.245 81.025 ;
        RECT 280.860 80.980 281.150 81.025 ;
        RECT 282.315 81.025 294.965 81.165 ;
        RECT 266.215 80.825 266.355 80.965 ;
        RECT 260.650 80.685 264.515 80.825 ;
        RECT 256.020 80.345 257.245 80.485 ;
        RECT 256.020 80.300 256.310 80.345 ;
        RECT 256.925 80.285 257.245 80.345 ;
        RECT 257.400 80.300 257.690 80.530 ;
        RECT 257.845 80.485 258.165 80.545 ;
        RECT 258.855 80.530 258.995 80.685 ;
        RECT 260.145 80.625 260.465 80.685 ;
        RECT 257.845 80.345 258.360 80.485 ;
        RECT 257.845 80.285 258.165 80.345 ;
        RECT 258.780 80.300 259.070 80.530 ;
        RECT 259.225 80.285 259.545 80.545 ;
        RECT 259.725 80.300 260.015 80.530 ;
        RECT 260.235 80.485 260.375 80.625 ;
        RECT 261.770 80.485 262.060 80.530 ;
        RECT 260.235 80.345 262.060 80.485 ;
        RECT 261.770 80.300 262.060 80.345 ;
        RECT 244.505 79.945 244.825 80.205 ;
        RECT 256.465 80.145 256.785 80.205 ;
        RECT 259.800 80.145 259.940 80.300 ;
        RECT 262.445 80.285 262.765 80.545 ;
        RECT 262.920 80.485 263.210 80.530 ;
        RECT 262.920 80.345 263.595 80.485 ;
        RECT 262.920 80.300 263.210 80.345 ;
        RECT 256.465 80.005 259.940 80.145 ;
        RECT 263.455 80.145 263.595 80.345 ;
        RECT 263.825 80.285 264.145 80.545 ;
        RECT 264.375 80.530 264.515 80.685 ;
        RECT 265.755 80.685 266.355 80.825 ;
        RECT 265.755 80.530 265.895 80.685 ;
        RECT 268.425 80.625 268.745 80.885 ;
        RECT 282.315 80.825 282.455 81.025 ;
        RECT 292.345 80.965 292.665 81.025 ;
        RECT 294.645 80.965 294.965 81.025 ;
        RECT 297.520 81.165 297.810 81.210 ;
        RECT 300.640 81.165 300.930 81.210 ;
        RECT 302.530 81.165 302.820 81.210 ;
        RECT 297.520 81.025 302.820 81.165 ;
        RECT 297.520 80.980 297.810 81.025 ;
        RECT 300.640 80.980 300.930 81.025 ;
        RECT 302.530 80.980 302.820 81.025 ;
        RECT 279.555 80.685 282.455 80.825 ;
        RECT 283.145 80.825 283.465 80.885 ;
        RECT 283.620 80.825 283.910 80.870 ;
        RECT 287.760 80.825 288.050 80.870 ;
        RECT 283.145 80.685 288.050 80.825 ;
        RECT 264.300 80.300 264.590 80.530 ;
        RECT 265.680 80.300 265.970 80.530 ;
        RECT 266.125 80.285 266.445 80.545 ;
        RECT 266.600 80.485 266.890 80.530 ;
        RECT 267.045 80.485 267.365 80.545 ;
        RECT 266.600 80.345 267.365 80.485 ;
        RECT 266.600 80.300 266.890 80.345 ;
        RECT 266.675 80.145 266.815 80.300 ;
        RECT 267.045 80.285 267.365 80.345 ;
        RECT 267.505 80.285 267.825 80.545 ;
        RECT 267.980 80.300 268.270 80.530 ;
        RECT 263.455 80.005 266.815 80.145 ;
        RECT 256.465 79.945 256.785 80.005 ;
        RECT 231.625 79.805 231.945 79.865 ;
        RECT 229.850 79.665 231.945 79.805 ;
        RECT 228.405 79.605 228.725 79.665 ;
        RECT 228.880 79.620 229.170 79.665 ;
        RECT 231.625 79.605 231.945 79.665 ;
        RECT 232.545 79.605 232.865 79.865 ;
        RECT 242.220 79.805 242.510 79.850 ;
        RECT 245.425 79.805 245.745 79.865 ;
        RECT 242.220 79.665 245.745 79.805 ;
        RECT 242.220 79.620 242.510 79.665 ;
        RECT 245.425 79.605 245.745 79.665 ;
        RECT 245.900 79.805 246.190 79.850 ;
        RECT 246.345 79.805 246.665 79.865 ;
        RECT 247.725 79.850 248.045 79.865 ;
        RECT 247.695 79.805 248.045 79.850 ;
        RECT 250.485 79.805 250.805 79.865 ;
        RECT 245.900 79.665 246.665 79.805 ;
        RECT 247.530 79.665 250.805 79.805 ;
        RECT 245.900 79.620 246.190 79.665 ;
        RECT 246.345 79.605 246.665 79.665 ;
        RECT 247.695 79.620 248.045 79.665 ;
        RECT 247.725 79.605 248.045 79.620 ;
        RECT 250.485 79.605 250.805 79.665 ;
        RECT 260.620 79.805 260.910 79.850 ;
        RECT 268.055 79.805 268.195 80.300 ;
        RECT 269.345 80.285 269.665 80.545 ;
        RECT 268.885 80.145 269.205 80.205 ;
        RECT 279.555 80.145 279.695 80.685 ;
        RECT 283.145 80.625 283.465 80.685 ;
        RECT 283.620 80.640 283.910 80.685 ;
        RECT 287.760 80.640 288.050 80.685 ;
        RECT 290.965 80.625 291.285 80.885 ;
        RECT 296.025 80.825 296.345 80.885 ;
        RECT 303.400 80.825 303.690 80.870 ;
        RECT 296.025 80.685 303.690 80.825 ;
        RECT 296.025 80.625 296.345 80.685 ;
        RECT 303.400 80.640 303.690 80.685 ;
        RECT 280.385 80.485 280.705 80.545 ;
        RECT 287.300 80.485 287.590 80.530 ;
        RECT 280.385 80.345 287.590 80.485 ;
        RECT 280.385 80.285 280.705 80.345 ;
        RECT 287.300 80.300 287.590 80.345 ;
        RECT 291.885 80.285 292.205 80.545 ;
        RECT 268.885 80.005 279.695 80.145 ;
        RECT 283.160 80.145 283.450 80.190 ;
        RECT 283.605 80.145 283.925 80.205 ;
        RECT 296.440 80.190 296.730 80.505 ;
        RECT 297.520 80.485 297.810 80.530 ;
        RECT 301.100 80.485 301.390 80.530 ;
        RECT 302.935 80.485 303.225 80.530 ;
        RECT 297.520 80.345 303.225 80.485 ;
        RECT 297.520 80.300 297.810 80.345 ;
        RECT 301.100 80.300 301.390 80.345 ;
        RECT 302.935 80.300 303.225 80.345 ;
        RECT 283.160 80.005 283.925 80.145 ;
        RECT 268.885 79.945 269.205 80.005 ;
        RECT 283.160 79.960 283.450 80.005 ;
        RECT 283.605 79.945 283.925 80.005 ;
        RECT 296.140 80.145 296.730 80.190 ;
        RECT 299.380 80.145 300.030 80.190 ;
        RECT 302.020 80.145 302.310 80.190 ;
        RECT 304.305 80.145 304.625 80.205 ;
        RECT 296.140 80.005 300.855 80.145 ;
        RECT 296.140 79.960 296.430 80.005 ;
        RECT 299.380 79.960 300.030 80.005 ;
        RECT 260.620 79.665 268.195 79.805 ;
        RECT 260.620 79.620 260.910 79.665 ;
        RECT 270.265 79.605 270.585 79.865 ;
        RECT 281.305 79.805 281.625 79.865 ;
        RECT 282.700 79.805 282.990 79.850 ;
        RECT 281.305 79.665 282.990 79.805 ;
        RECT 281.305 79.605 281.625 79.665 ;
        RECT 282.700 79.620 282.990 79.665 ;
        RECT 284.985 79.605 285.305 79.865 ;
        RECT 286.840 79.805 287.130 79.850 ;
        RECT 289.125 79.805 289.445 79.865 ;
        RECT 286.840 79.665 289.445 79.805 ;
        RECT 286.840 79.620 287.130 79.665 ;
        RECT 289.125 79.605 289.445 79.665 ;
        RECT 292.345 79.605 292.665 79.865 ;
        RECT 294.185 79.605 294.505 79.865 ;
        RECT 300.715 79.805 300.855 80.005 ;
        RECT 302.020 80.005 304.625 80.145 ;
        RECT 302.020 79.960 302.310 80.005 ;
        RECT 304.305 79.945 304.625 80.005 ;
        RECT 302.465 79.805 302.785 79.865 ;
        RECT 300.715 79.665 302.785 79.805 ;
        RECT 302.465 79.605 302.785 79.665 ;
        RECT 162.095 78.985 311.135 79.465 ;
        RECT 178.740 78.785 179.030 78.830 ;
        RECT 181.960 78.785 182.250 78.830 ;
        RECT 182.865 78.785 183.185 78.845 ;
        RECT 178.740 78.645 183.185 78.785 ;
        RECT 178.740 78.600 179.030 78.645 ;
        RECT 181.960 78.600 182.250 78.645 ;
        RECT 182.865 78.585 183.185 78.645 ;
        RECT 183.785 78.785 184.105 78.845 ;
        RECT 193.905 78.785 194.225 78.845 ;
        RECT 183.785 78.645 194.225 78.785 ;
        RECT 183.785 78.585 184.105 78.645 ;
        RECT 193.905 78.585 194.225 78.645 ;
        RECT 195.745 78.785 196.065 78.845 ;
        RECT 200.345 78.785 200.665 78.845 ;
        RECT 215.065 78.785 215.385 78.845 ;
        RECT 220.125 78.785 220.445 78.845 ;
        RECT 195.745 78.645 200.665 78.785 ;
        RECT 195.745 78.585 196.065 78.645 ;
        RECT 173.660 78.445 174.310 78.490 ;
        RECT 177.260 78.445 177.550 78.490 ;
        RECT 173.660 78.305 177.550 78.445 ;
        RECT 173.660 78.260 174.310 78.305 ;
        RECT 176.960 78.260 177.550 78.305 ;
        RECT 180.565 78.445 180.885 78.505 ;
        RECT 189.320 78.445 189.610 78.490 ;
        RECT 180.565 78.305 189.610 78.445 ;
        RECT 176.960 78.165 177.250 78.260 ;
        RECT 180.565 78.245 180.885 78.305 ;
        RECT 189.320 78.260 189.610 78.305 ;
        RECT 193.445 78.245 193.765 78.505 ;
        RECT 195.285 78.445 195.605 78.505 ;
        RECT 198.595 78.445 198.735 78.645 ;
        RECT 200.345 78.585 200.665 78.645 ;
        RECT 204.575 78.645 220.445 78.785 ;
        RECT 204.575 78.490 204.715 78.645 ;
        RECT 215.065 78.585 215.385 78.645 ;
        RECT 220.125 78.585 220.445 78.645 ;
        RECT 220.585 78.785 220.905 78.845 ;
        RECT 227.945 78.785 228.265 78.845 ;
        RECT 220.585 78.645 228.265 78.785 ;
        RECT 220.585 78.585 220.905 78.645 ;
        RECT 227.945 78.585 228.265 78.645 ;
        RECT 228.865 78.830 229.185 78.845 ;
        RECT 228.865 78.785 229.215 78.830 ;
        RECT 260.605 78.785 260.925 78.845 ;
        RECT 261.080 78.785 261.370 78.830 ;
        RECT 228.865 78.645 229.380 78.785 ;
        RECT 243.675 78.645 259.455 78.785 ;
        RECT 228.865 78.600 229.215 78.645 ;
        RECT 228.865 78.585 229.185 78.600 ;
        RECT 204.500 78.445 204.790 78.490 ;
        RECT 195.285 78.305 197.355 78.445 ;
        RECT 195.285 78.245 195.605 78.305 ;
        RECT 197.215 78.165 197.355 78.305 ;
        RECT 198.135 78.305 198.735 78.445 ;
        RECT 199.975 78.305 204.790 78.445 ;
        RECT 165.845 78.105 166.165 78.165 ;
        RECT 170.000 78.105 170.290 78.150 ;
        RECT 165.845 77.965 170.290 78.105 ;
        RECT 165.845 77.905 166.165 77.965 ;
        RECT 170.000 77.920 170.290 77.965 ;
        RECT 170.465 78.105 170.755 78.150 ;
        RECT 172.300 78.105 172.590 78.150 ;
        RECT 175.880 78.105 176.170 78.150 ;
        RECT 170.465 77.965 176.170 78.105 ;
        RECT 170.465 77.920 170.755 77.965 ;
        RECT 172.300 77.920 172.590 77.965 ;
        RECT 175.880 77.920 176.170 77.965 ;
        RECT 176.885 77.945 177.250 78.165 ;
        RECT 179.645 78.105 179.965 78.165 ;
        RECT 179.645 77.965 180.335 78.105 ;
        RECT 176.885 77.905 177.205 77.945 ;
        RECT 179.645 77.905 179.965 77.965 ;
        RECT 171.380 77.765 171.670 77.810 ;
        RECT 171.380 77.625 179.875 77.765 ;
        RECT 171.380 77.580 171.670 77.625 ;
        RECT 179.735 77.470 179.875 77.625 ;
        RECT 170.870 77.425 171.160 77.470 ;
        RECT 172.760 77.425 173.050 77.470 ;
        RECT 175.880 77.425 176.170 77.470 ;
        RECT 170.870 77.285 176.170 77.425 ;
        RECT 170.870 77.240 171.160 77.285 ;
        RECT 172.760 77.240 173.050 77.285 ;
        RECT 175.880 77.240 176.170 77.285 ;
        RECT 179.660 77.240 179.950 77.470 ;
        RECT 180.195 77.425 180.335 77.965 ;
        RECT 181.485 77.905 181.805 78.165 ;
        RECT 185.640 78.105 185.930 78.150 ;
        RECT 187.005 78.105 187.325 78.165 ;
        RECT 185.640 77.965 187.325 78.105 ;
        RECT 185.640 77.920 185.930 77.965 ;
        RECT 187.005 77.905 187.325 77.965 ;
        RECT 187.480 78.105 187.770 78.150 ;
        RECT 187.925 78.105 188.245 78.165 ;
        RECT 193.920 78.105 194.210 78.150 ;
        RECT 187.480 77.965 188.245 78.105 ;
        RECT 187.480 77.920 187.770 77.965 ;
        RECT 187.925 77.905 188.245 77.965 ;
        RECT 189.395 77.965 196.435 78.105 ;
        RECT 189.395 77.825 189.535 77.965 ;
        RECT 193.920 77.920 194.210 77.965 ;
        RECT 182.880 77.580 183.170 77.810 ;
        RECT 182.955 77.425 183.095 77.580 ;
        RECT 184.705 77.565 185.025 77.825 ;
        RECT 189.305 77.565 189.625 77.825 ;
        RECT 194.365 77.565 194.685 77.825 ;
        RECT 196.295 77.765 196.435 77.965 ;
        RECT 196.665 77.905 196.985 78.165 ;
        RECT 197.125 78.105 197.445 78.165 ;
        RECT 198.135 78.150 198.275 78.305 ;
        RECT 197.600 78.105 197.890 78.150 ;
        RECT 197.125 77.965 197.890 78.105 ;
        RECT 197.125 77.905 197.445 77.965 ;
        RECT 197.600 77.920 197.890 77.965 ;
        RECT 198.060 77.920 198.350 78.150 ;
        RECT 198.520 78.105 198.810 78.150 ;
        RECT 198.965 78.105 199.285 78.165 ;
        RECT 198.520 77.965 199.285 78.105 ;
        RECT 198.520 77.920 198.810 77.965 ;
        RECT 198.965 77.905 199.285 77.965 ;
        RECT 199.975 77.765 200.115 78.305 ;
        RECT 204.500 78.260 204.790 78.305 ;
        RECT 204.945 78.445 205.265 78.505 ;
        RECT 206.385 78.445 206.675 78.490 ;
        RECT 204.945 78.305 206.675 78.445 ;
        RECT 204.945 78.245 205.265 78.305 ;
        RECT 206.385 78.260 206.675 78.305 ;
        RECT 207.245 78.445 207.565 78.505 ;
        RECT 228.405 78.445 228.725 78.505 ;
        RECT 233.925 78.445 234.245 78.505 ;
        RECT 243.675 78.490 243.815 78.645 ;
        RECT 243.600 78.445 243.890 78.490 ;
        RECT 207.245 78.305 224.955 78.445 ;
        RECT 207.245 78.245 207.565 78.305 ;
        RECT 202.185 78.105 202.505 78.165 ;
        RECT 210.005 78.105 210.325 78.165 ;
        RECT 202.185 77.965 210.325 78.105 ;
        RECT 202.185 77.905 202.505 77.965 ;
        RECT 210.005 77.905 210.325 77.965 ;
        RECT 210.940 77.920 211.230 78.150 ;
        RECT 211.860 78.105 212.150 78.150 ;
        RECT 212.305 78.105 212.625 78.165 ;
        RECT 224.815 78.150 224.955 78.305 ;
        RECT 225.735 78.305 228.725 78.445 ;
        RECT 225.735 78.150 225.875 78.305 ;
        RECT 228.405 78.245 228.725 78.305 ;
        RECT 230.335 78.305 243.890 78.445 ;
        RECT 211.860 77.965 212.625 78.105 ;
        RECT 211.860 77.920 212.150 77.965 ;
        RECT 196.295 77.625 200.115 77.765 ;
        RECT 200.345 77.765 200.665 77.825 ;
        RECT 210.465 77.765 210.785 77.825 ;
        RECT 211.015 77.765 211.155 77.920 ;
        RECT 212.305 77.905 212.625 77.965 ;
        RECT 224.740 77.920 225.030 78.150 ;
        RECT 225.660 77.920 225.950 78.150 ;
        RECT 227.040 78.105 227.330 78.150 ;
        RECT 227.485 78.105 227.805 78.165 ;
        RECT 230.335 78.150 230.475 78.305 ;
        RECT 233.925 78.245 234.245 78.305 ;
        RECT 243.600 78.260 243.890 78.305 ;
        RECT 245.425 78.445 245.745 78.505 ;
        RECT 245.900 78.445 246.190 78.490 ;
        RECT 248.645 78.445 248.965 78.505 ;
        RECT 245.425 78.305 246.190 78.445 ;
        RECT 245.425 78.245 245.745 78.305 ;
        RECT 245.900 78.260 246.190 78.305 ;
        RECT 246.335 78.305 248.965 78.445 ;
        RECT 227.040 77.965 227.805 78.105 ;
        RECT 227.040 77.920 227.330 77.965 ;
        RECT 227.485 77.905 227.805 77.965 ;
        RECT 230.260 77.920 230.550 78.150 ;
        RECT 231.625 78.105 231.945 78.165 ;
        RECT 242.205 78.105 242.525 78.165 ;
        RECT 242.680 78.105 242.970 78.150 ;
        RECT 231.625 77.965 233.235 78.105 ;
        RECT 231.625 77.905 231.945 77.965 ;
        RECT 200.345 77.625 211.155 77.765 ;
        RECT 211.385 77.765 211.705 77.825 ;
        RECT 226.120 77.765 226.410 77.810 ;
        RECT 232.545 77.765 232.865 77.825 ;
        RECT 211.385 77.625 218.975 77.765 ;
        RECT 200.345 77.565 200.665 77.625 ;
        RECT 210.465 77.565 210.785 77.625 ;
        RECT 211.385 77.565 211.705 77.625 ;
        RECT 186.545 77.425 186.865 77.485 ;
        RECT 218.285 77.425 218.605 77.485 ;
        RECT 180.195 77.285 186.865 77.425 ;
        RECT 186.545 77.225 186.865 77.285 ;
        RECT 193.535 77.285 218.605 77.425 ;
        RECT 180.105 77.085 180.425 77.145 ;
        RECT 181.485 77.085 181.805 77.145 ;
        RECT 193.535 77.085 193.675 77.285 ;
        RECT 218.285 77.225 218.605 77.285 ;
        RECT 180.105 76.945 193.675 77.085 ;
        RECT 180.105 76.885 180.425 76.945 ;
        RECT 181.485 76.885 181.805 76.945 ;
        RECT 193.905 76.885 194.225 77.145 ;
        RECT 199.900 77.085 200.190 77.130 ;
        RECT 201.725 77.085 202.045 77.145 ;
        RECT 199.900 76.945 202.045 77.085 ;
        RECT 199.900 76.900 200.190 76.945 ;
        RECT 201.725 76.885 202.045 76.945 ;
        RECT 206.325 76.885 206.645 77.145 ;
        RECT 206.785 77.085 207.105 77.145 ;
        RECT 207.260 77.085 207.550 77.130 ;
        RECT 206.785 76.945 207.550 77.085 ;
        RECT 206.785 76.885 207.105 76.945 ;
        RECT 207.260 76.900 207.550 76.945 ;
        RECT 212.765 76.885 213.085 77.145 ;
        RECT 218.835 77.085 218.975 77.625 ;
        RECT 226.120 77.625 232.865 77.765 ;
        RECT 233.095 77.765 233.235 77.965 ;
        RECT 242.205 77.965 242.970 78.105 ;
        RECT 242.205 77.905 242.525 77.965 ;
        RECT 242.680 77.920 242.970 77.965 ;
        RECT 244.045 77.905 244.365 78.165 ;
        RECT 244.520 78.105 244.810 78.150 ;
        RECT 246.335 78.105 246.475 78.305 ;
        RECT 248.645 78.245 248.965 78.305 ;
        RECT 256.465 78.445 256.785 78.505 ;
        RECT 259.315 78.445 259.455 78.645 ;
        RECT 260.605 78.645 261.370 78.785 ;
        RECT 260.605 78.585 260.925 78.645 ;
        RECT 261.080 78.600 261.370 78.645 ;
        RECT 261.985 78.585 262.305 78.845 ;
        RECT 264.300 78.785 264.590 78.830 ;
        RECT 268.425 78.785 268.745 78.845 ;
        RECT 279.940 78.785 280.230 78.830 ;
        RECT 280.385 78.785 280.705 78.845 ;
        RECT 292.345 78.785 292.665 78.845 ;
        RECT 264.300 78.645 268.745 78.785 ;
        RECT 264.300 78.600 264.590 78.645 ;
        RECT 268.425 78.585 268.745 78.645 ;
        RECT 269.665 78.645 280.705 78.785 ;
        RECT 262.075 78.445 262.215 78.585 ;
        RECT 265.205 78.445 265.525 78.505 ;
        RECT 265.680 78.445 265.970 78.490 ;
        RECT 256.465 78.305 258.900 78.445 ;
        RECT 259.315 78.305 260.375 78.445 ;
        RECT 262.075 78.305 263.595 78.445 ;
        RECT 256.465 78.245 256.785 78.305 ;
        RECT 244.520 77.965 246.475 78.105 ;
        RECT 244.520 77.920 244.810 77.965 ;
        RECT 244.595 77.765 244.735 77.920 ;
        RECT 247.265 77.905 247.585 78.165 ;
        RECT 258.320 77.920 258.610 78.150 ;
        RECT 258.760 78.105 258.900 78.305 ;
        RECT 260.235 78.150 260.375 78.305 ;
        RECT 258.760 78.095 258.995 78.105 ;
        RECT 259.240 78.095 259.530 78.150 ;
        RECT 258.760 77.965 259.530 78.095 ;
        RECT 258.855 77.955 259.530 77.965 ;
        RECT 259.240 77.920 259.530 77.955 ;
        RECT 259.700 77.920 259.990 78.150 ;
        RECT 260.160 78.105 260.450 78.150 ;
        RECT 261.540 78.105 261.830 78.150 ;
        RECT 261.985 78.105 262.305 78.165 ;
        RECT 263.455 78.150 263.595 78.305 ;
        RECT 265.205 78.305 265.970 78.445 ;
        RECT 265.205 78.245 265.525 78.305 ;
        RECT 265.680 78.260 265.970 78.305 ;
        RECT 260.160 77.965 261.320 78.105 ;
        RECT 260.160 77.920 260.450 77.965 ;
        RECT 233.095 77.625 244.735 77.765 ;
        RECT 226.120 77.580 226.410 77.625 ;
        RECT 232.545 77.565 232.865 77.625 ;
        RECT 246.345 77.565 246.665 77.825 ;
        RECT 223.820 77.425 224.110 77.470 ;
        RECT 226.565 77.425 226.885 77.485 ;
        RECT 256.465 77.425 256.785 77.485 ;
        RECT 258.395 77.425 258.535 77.920 ;
        RECT 259.775 77.765 259.915 77.920 ;
        RECT 260.605 77.765 260.925 77.825 ;
        RECT 259.775 77.625 260.925 77.765 ;
        RECT 261.180 77.765 261.320 77.965 ;
        RECT 261.540 77.965 262.305 78.105 ;
        RECT 261.540 77.920 261.830 77.965 ;
        RECT 261.985 77.905 262.305 77.965 ;
        RECT 262.460 77.920 262.750 78.150 ;
        RECT 262.920 77.920 263.210 78.150 ;
        RECT 263.380 78.105 263.670 78.150 ;
        RECT 266.600 78.105 266.890 78.150 ;
        RECT 263.380 77.965 266.890 78.105 ;
        RECT 263.380 77.920 263.670 77.965 ;
        RECT 266.600 77.920 266.890 77.965 ;
        RECT 267.965 78.105 268.285 78.165 ;
        RECT 269.665 78.105 269.805 78.645 ;
        RECT 279.940 78.600 280.230 78.645 ;
        RECT 280.385 78.585 280.705 78.645 ;
        RECT 280.935 78.645 292.665 78.785 ;
        RECT 267.965 77.965 269.805 78.105 ;
        RECT 262.535 77.765 262.675 77.920 ;
        RECT 261.180 77.625 262.675 77.765 ;
        RECT 260.605 77.565 260.925 77.625 ;
        RECT 223.820 77.285 226.885 77.425 ;
        RECT 223.820 77.240 224.110 77.285 ;
        RECT 226.565 77.225 226.885 77.285 ;
        RECT 227.575 77.285 258.535 77.425 ;
        RECT 262.995 77.425 263.135 77.920 ;
        RECT 267.965 77.905 268.285 77.965 ;
        RECT 264.285 77.765 264.605 77.825 ;
        RECT 267.520 77.765 267.810 77.810 ;
        RECT 272.565 77.765 272.885 77.825 ;
        RECT 280.935 77.765 281.075 78.645 ;
        RECT 292.345 78.585 292.665 78.645 ;
        RECT 306.605 78.585 306.925 78.845 ;
        RECT 281.420 78.445 281.710 78.490 ;
        RECT 284.065 78.445 284.385 78.505 ;
        RECT 284.660 78.445 285.310 78.490 ;
        RECT 281.420 78.305 285.310 78.445 ;
        RECT 281.420 78.260 282.010 78.305 ;
        RECT 281.720 77.945 282.010 78.260 ;
        RECT 284.065 78.245 284.385 78.305 ;
        RECT 284.660 78.260 285.310 78.305 ;
        RECT 287.285 78.445 287.605 78.505 ;
        RECT 289.585 78.445 289.905 78.505 ;
        RECT 291.440 78.445 291.730 78.490 ;
        RECT 287.285 78.305 291.730 78.445 ;
        RECT 287.285 78.245 287.605 78.305 ;
        RECT 289.585 78.245 289.905 78.305 ;
        RECT 291.440 78.260 291.730 78.305 ;
        RECT 301.540 78.445 302.190 78.490 ;
        RECT 302.465 78.445 302.785 78.505 ;
        RECT 305.140 78.445 305.430 78.490 ;
        RECT 301.540 78.305 305.430 78.445 ;
        RECT 301.540 78.260 302.190 78.305 ;
        RECT 302.465 78.245 302.785 78.305 ;
        RECT 304.840 78.260 305.430 78.305 ;
        RECT 282.800 78.105 283.090 78.150 ;
        RECT 286.380 78.105 286.670 78.150 ;
        RECT 288.215 78.105 288.505 78.150 ;
        RECT 282.800 77.965 288.505 78.105 ;
        RECT 282.800 77.920 283.090 77.965 ;
        RECT 286.380 77.920 286.670 77.965 ;
        RECT 288.215 77.920 288.505 77.965 ;
        RECT 288.680 78.105 288.970 78.150 ;
        RECT 290.505 78.105 290.825 78.165 ;
        RECT 296.025 78.105 296.345 78.165 ;
        RECT 297.880 78.105 298.170 78.150 ;
        RECT 288.680 77.965 298.170 78.105 ;
        RECT 288.680 77.920 288.970 77.965 ;
        RECT 290.505 77.905 290.825 77.965 ;
        RECT 296.025 77.905 296.345 77.965 ;
        RECT 297.880 77.920 298.170 77.965 ;
        RECT 298.345 78.105 298.635 78.150 ;
        RECT 300.180 78.105 300.470 78.150 ;
        RECT 303.760 78.105 304.050 78.150 ;
        RECT 298.345 77.965 304.050 78.105 ;
        RECT 298.345 77.920 298.635 77.965 ;
        RECT 300.180 77.920 300.470 77.965 ;
        RECT 303.760 77.920 304.050 77.965 ;
        RECT 304.840 77.945 305.130 78.260 ;
        RECT 264.285 77.625 281.075 77.765 ;
        RECT 284.985 77.765 285.305 77.825 ;
        RECT 287.300 77.765 287.590 77.810 ;
        RECT 284.985 77.625 287.590 77.765 ;
        RECT 264.285 77.565 264.605 77.625 ;
        RECT 267.520 77.580 267.810 77.625 ;
        RECT 272.565 77.565 272.885 77.625 ;
        RECT 284.985 77.565 285.305 77.625 ;
        RECT 287.300 77.580 287.590 77.625 ;
        RECT 295.105 77.565 295.425 77.825 ;
        RECT 299.260 77.765 299.550 77.810 ;
        RECT 299.260 77.625 304.995 77.765 ;
        RECT 299.260 77.580 299.550 77.625 ;
        RECT 304.855 77.485 304.995 77.625 ;
        RECT 268.425 77.425 268.745 77.485 ;
        RECT 282.800 77.425 283.090 77.470 ;
        RECT 285.920 77.425 286.210 77.470 ;
        RECT 287.810 77.425 288.100 77.470 ;
        RECT 262.995 77.285 268.745 77.425 ;
        RECT 227.575 77.085 227.715 77.285 ;
        RECT 256.465 77.225 256.785 77.285 ;
        RECT 268.425 77.225 268.745 77.285 ;
        RECT 269.435 77.285 282.455 77.425 ;
        RECT 218.835 76.945 227.715 77.085 ;
        RECT 228.880 77.085 229.170 77.130 ;
        RECT 229.325 77.085 229.645 77.145 ;
        RECT 228.880 76.945 229.645 77.085 ;
        RECT 228.880 76.900 229.170 76.945 ;
        RECT 229.325 76.885 229.645 76.945 ;
        RECT 245.440 77.085 245.730 77.130 ;
        RECT 245.900 77.085 246.190 77.130 ;
        RECT 245.440 76.945 246.190 77.085 ;
        RECT 245.440 76.900 245.730 76.945 ;
        RECT 245.900 76.900 246.190 76.945 ;
        RECT 248.185 76.885 248.505 77.145 ;
        RECT 258.305 77.085 258.625 77.145 ;
        RECT 259.685 77.085 260.005 77.145 ;
        RECT 258.305 76.945 260.005 77.085 ;
        RECT 258.305 76.885 258.625 76.945 ;
        RECT 259.685 76.885 260.005 76.945 ;
        RECT 261.985 77.085 262.305 77.145 ;
        RECT 269.435 77.085 269.575 77.285 ;
        RECT 261.985 76.945 269.575 77.085 ;
        RECT 282.315 77.085 282.455 77.285 ;
        RECT 282.800 77.285 288.100 77.425 ;
        RECT 282.800 77.240 283.090 77.285 ;
        RECT 285.920 77.240 286.210 77.285 ;
        RECT 287.810 77.240 288.100 77.285 ;
        RECT 298.750 77.425 299.040 77.470 ;
        RECT 300.640 77.425 300.930 77.470 ;
        RECT 303.760 77.425 304.050 77.470 ;
        RECT 298.750 77.285 304.050 77.425 ;
        RECT 298.750 77.240 299.040 77.285 ;
        RECT 300.640 77.240 300.930 77.285 ;
        RECT 303.760 77.240 304.050 77.285 ;
        RECT 304.765 77.225 305.085 77.485 ;
        RECT 288.665 77.085 288.985 77.145 ;
        RECT 282.315 76.945 288.985 77.085 ;
        RECT 261.985 76.885 262.305 76.945 ;
        RECT 288.665 76.885 288.985 76.945 ;
        RECT 294.645 77.085 294.965 77.145 ;
        RECT 302.925 77.085 303.245 77.145 ;
        RECT 294.645 76.945 303.245 77.085 ;
        RECT 294.645 76.885 294.965 76.945 ;
        RECT 302.925 76.885 303.245 76.945 ;
        RECT 162.095 76.265 311.135 76.745 ;
        RECT 167.175 76.065 167.465 76.110 ;
        RECT 175.520 76.065 175.810 76.110 ;
        RECT 167.175 75.925 175.810 76.065 ;
        RECT 167.175 75.880 167.465 75.925 ;
        RECT 175.520 75.880 175.810 75.925 ;
        RECT 176.885 76.065 177.205 76.125 ;
        RECT 189.780 76.065 190.070 76.110 ;
        RECT 190.685 76.065 191.005 76.125 ;
        RECT 199.425 76.065 199.745 76.125 ;
        RECT 176.885 75.925 188.615 76.065 ;
        RECT 176.885 75.865 177.205 75.925 ;
        RECT 166.730 75.725 167.020 75.770 ;
        RECT 168.620 75.725 168.910 75.770 ;
        RECT 171.740 75.725 172.030 75.770 ;
        RECT 166.730 75.585 172.030 75.725 ;
        RECT 166.730 75.540 167.020 75.585 ;
        RECT 168.620 75.540 168.910 75.585 ;
        RECT 171.740 75.540 172.030 75.585 ;
        RECT 181.910 75.725 182.200 75.770 ;
        RECT 183.800 75.725 184.090 75.770 ;
        RECT 186.920 75.725 187.210 75.770 ;
        RECT 181.910 75.585 187.210 75.725 ;
        RECT 181.910 75.540 182.200 75.585 ;
        RECT 183.800 75.540 184.090 75.585 ;
        RECT 186.920 75.540 187.210 75.585 ;
        RECT 165.860 75.385 166.150 75.430 ;
        RECT 173.205 75.385 173.525 75.445 ;
        RECT 165.860 75.245 173.525 75.385 ;
        RECT 165.860 75.200 166.150 75.245 ;
        RECT 173.205 75.185 173.525 75.245 ;
        RECT 174.600 75.385 174.890 75.430 ;
        RECT 178.740 75.385 179.030 75.430 ;
        RECT 179.645 75.385 179.965 75.445 ;
        RECT 174.600 75.245 178.035 75.385 ;
        RECT 174.600 75.200 174.890 75.245 ;
        RECT 166.325 75.045 166.615 75.090 ;
        RECT 168.160 75.045 168.450 75.090 ;
        RECT 171.740 75.045 172.030 75.090 ;
        RECT 166.325 74.905 172.030 75.045 ;
        RECT 166.325 74.860 166.615 74.905 ;
        RECT 168.160 74.860 168.450 74.905 ;
        RECT 171.740 74.860 172.030 74.905 ;
        RECT 172.820 74.750 173.110 75.065 ;
        RECT 169.520 74.705 170.170 74.750 ;
        RECT 172.820 74.705 173.410 74.750 ;
        RECT 173.665 74.705 173.985 74.765 ;
        RECT 176.885 74.705 177.205 74.765 ;
        RECT 177.895 74.750 178.035 75.245 ;
        RECT 178.740 75.245 179.965 75.385 ;
        RECT 178.740 75.200 179.030 75.245 ;
        RECT 179.645 75.185 179.965 75.245 ;
        RECT 180.565 75.385 180.885 75.445 ;
        RECT 181.040 75.385 181.330 75.430 ;
        RECT 182.865 75.385 183.185 75.445 ;
        RECT 180.565 75.245 183.185 75.385 ;
        RECT 180.565 75.185 180.885 75.245 ;
        RECT 181.040 75.200 181.330 75.245 ;
        RECT 182.865 75.185 183.185 75.245 ;
        RECT 181.505 75.045 181.795 75.090 ;
        RECT 183.340 75.045 183.630 75.090 ;
        RECT 186.920 75.045 187.210 75.090 ;
        RECT 181.505 74.905 187.210 75.045 ;
        RECT 181.505 74.860 181.795 74.905 ;
        RECT 183.340 74.860 183.630 74.905 ;
        RECT 186.920 74.860 187.210 74.905 ;
        RECT 169.520 74.565 177.205 74.705 ;
        RECT 169.520 74.520 170.170 74.565 ;
        RECT 173.120 74.520 173.410 74.565 ;
        RECT 173.665 74.505 173.985 74.565 ;
        RECT 176.885 74.505 177.205 74.565 ;
        RECT 177.820 74.705 178.110 74.750 ;
        RECT 181.025 74.705 181.345 74.765 ;
        RECT 188.000 74.750 188.290 75.065 ;
        RECT 188.475 74.750 188.615 75.925 ;
        RECT 189.780 75.925 199.745 76.065 ;
        RECT 189.780 75.880 190.070 75.925 ;
        RECT 190.685 75.865 191.005 75.925 ;
        RECT 199.425 75.865 199.745 75.925 ;
        RECT 200.345 76.065 200.665 76.125 ;
        RECT 202.185 76.065 202.505 76.125 ;
        RECT 212.305 76.065 212.625 76.125 ;
        RECT 221.965 76.065 222.285 76.125 ;
        RECT 224.280 76.065 224.570 76.110 ;
        RECT 200.345 75.925 202.505 76.065 ;
        RECT 200.345 75.865 200.665 75.925 ;
        RECT 202.185 75.865 202.505 75.925 ;
        RECT 202.735 75.925 224.570 76.065 ;
        RECT 192.490 75.725 192.780 75.770 ;
        RECT 194.380 75.725 194.670 75.770 ;
        RECT 197.500 75.725 197.790 75.770 ;
        RECT 192.490 75.585 197.790 75.725 ;
        RECT 192.490 75.540 192.780 75.585 ;
        RECT 194.380 75.540 194.670 75.585 ;
        RECT 197.500 75.540 197.790 75.585 ;
        RECT 191.605 75.185 191.925 75.445 ;
        RECT 202.735 75.090 202.875 75.925 ;
        RECT 212.305 75.865 212.625 75.925 ;
        RECT 221.965 75.865 222.285 75.925 ;
        RECT 224.280 75.880 224.570 75.925 ;
        RECT 243.585 76.065 243.905 76.125 ;
        RECT 258.305 76.065 258.625 76.125 ;
        RECT 264.285 76.065 264.605 76.125 ;
        RECT 243.585 75.925 256.005 76.065 ;
        RECT 243.585 75.865 243.905 75.925 ;
        RECT 205.405 75.725 205.725 75.785 ;
        RECT 207.260 75.725 207.550 75.770 ;
        RECT 205.405 75.585 207.550 75.725 ;
        RECT 205.405 75.525 205.725 75.585 ;
        RECT 207.260 75.540 207.550 75.585 ;
        RECT 210.120 75.725 210.410 75.770 ;
        RECT 213.240 75.725 213.530 75.770 ;
        RECT 215.130 75.725 215.420 75.770 ;
        RECT 210.120 75.585 215.420 75.725 ;
        RECT 210.120 75.540 210.410 75.585 ;
        RECT 213.240 75.540 213.530 75.585 ;
        RECT 215.130 75.540 215.420 75.585 ;
        RECT 216.460 75.725 216.750 75.770 ;
        RECT 216.905 75.725 217.225 75.785 ;
        RECT 216.460 75.585 217.225 75.725 ;
        RECT 216.460 75.540 216.750 75.585 ;
        RECT 192.085 75.045 192.375 75.090 ;
        RECT 193.920 75.045 194.210 75.090 ;
        RECT 197.500 75.045 197.790 75.090 ;
        RECT 192.085 74.905 197.790 75.045 ;
        RECT 192.085 74.860 192.375 74.905 ;
        RECT 193.920 74.860 194.210 74.905 ;
        RECT 197.500 74.860 197.790 74.905 ;
        RECT 177.820 74.565 181.345 74.705 ;
        RECT 177.820 74.520 178.110 74.565 ;
        RECT 181.025 74.505 181.345 74.565 ;
        RECT 182.420 74.520 182.710 74.750 ;
        RECT 184.700 74.705 185.350 74.750 ;
        RECT 188.000 74.705 188.615 74.750 ;
        RECT 193.000 74.705 193.290 74.750 ;
        RECT 194.365 74.705 194.685 74.765 ;
        RECT 198.580 74.750 198.870 75.065 ;
        RECT 202.660 74.860 202.950 75.090 ;
        RECT 195.280 74.705 195.930 74.750 ;
        RECT 198.580 74.705 199.170 74.750 ;
        RECT 184.700 74.565 192.755 74.705 ;
        RECT 184.700 74.520 185.350 74.565 ;
        RECT 188.300 74.520 188.590 74.565 ;
        RECT 177.345 74.165 177.665 74.425 ;
        RECT 182.495 74.365 182.635 74.520 ;
        RECT 192.615 74.425 192.755 74.565 ;
        RECT 193.000 74.565 194.685 74.705 ;
        RECT 193.000 74.520 193.290 74.565 ;
        RECT 194.365 74.505 194.685 74.565 ;
        RECT 194.915 74.565 199.170 74.705 ;
        RECT 188.845 74.365 189.165 74.425 ;
        RECT 182.495 74.225 189.165 74.365 ;
        RECT 188.845 74.165 189.165 74.225 ;
        RECT 192.525 74.365 192.845 74.425 ;
        RECT 194.915 74.365 195.055 74.565 ;
        RECT 195.280 74.520 195.930 74.565 ;
        RECT 198.880 74.520 199.170 74.565 ;
        RECT 201.740 74.365 202.030 74.410 ;
        RECT 192.525 74.225 202.030 74.365 ;
        RECT 207.335 74.365 207.475 75.540 ;
        RECT 216.905 75.525 217.225 75.585 ;
        RECT 218.745 75.725 219.065 75.785 ;
        RECT 248.185 75.725 248.505 75.785 ;
        RECT 218.745 75.585 248.505 75.725 ;
        RECT 255.865 75.725 256.005 75.925 ;
        RECT 258.305 75.925 264.605 76.065 ;
        RECT 258.305 75.865 258.625 75.925 ;
        RECT 264.285 75.865 264.605 75.925 ;
        RECT 292.345 76.065 292.665 76.125 ;
        RECT 303.400 76.065 303.690 76.110 ;
        RECT 292.345 75.925 303.690 76.065 ;
        RECT 292.345 75.865 292.665 75.925 ;
        RECT 303.400 75.880 303.690 75.925 ;
        RECT 304.305 75.865 304.625 76.125 ;
        RECT 262.445 75.725 262.765 75.785 ;
        RECT 263.365 75.725 263.685 75.785 ;
        RECT 255.865 75.585 262.215 75.725 ;
        RECT 218.745 75.525 219.065 75.585 ;
        RECT 248.185 75.525 248.505 75.585 ;
        RECT 211.845 75.385 212.165 75.445 ;
        RECT 216.000 75.385 216.290 75.430 ;
        RECT 211.845 75.245 216.290 75.385 ;
        RECT 211.845 75.185 212.165 75.245 ;
        RECT 216.000 75.200 216.290 75.245 ;
        RECT 217.825 75.385 218.145 75.445 ;
        RECT 219.220 75.385 219.510 75.430 ;
        RECT 217.825 75.245 219.510 75.385 ;
        RECT 209.040 74.750 209.330 75.065 ;
        RECT 210.120 75.045 210.410 75.090 ;
        RECT 213.700 75.045 213.990 75.090 ;
        RECT 215.535 75.045 215.825 75.090 ;
        RECT 210.120 74.905 215.825 75.045 ;
        RECT 216.075 75.045 216.215 75.200 ;
        RECT 217.825 75.185 218.145 75.245 ;
        RECT 219.220 75.200 219.510 75.245 ;
        RECT 227.945 75.385 228.265 75.445 ;
        RECT 261.065 75.385 261.385 75.445 ;
        RECT 227.945 75.245 261.385 75.385 ;
        RECT 227.945 75.185 228.265 75.245 ;
        RECT 225.200 75.045 225.490 75.090 ;
        RECT 238.525 75.045 238.845 75.105 ;
        RECT 216.075 74.905 219.435 75.045 ;
        RECT 210.120 74.860 210.410 74.905 ;
        RECT 213.700 74.860 213.990 74.905 ;
        RECT 215.535 74.860 215.825 74.905 ;
        RECT 219.295 74.765 219.435 74.905 ;
        RECT 225.200 74.905 238.845 75.045 ;
        RECT 225.200 74.860 225.490 74.905 ;
        RECT 238.525 74.845 238.845 74.905 ;
        RECT 244.965 75.045 245.285 75.105 ;
        RECT 247.725 75.045 248.045 75.105 ;
        RECT 244.965 74.905 248.045 75.045 ;
        RECT 244.965 74.845 245.285 74.905 ;
        RECT 247.725 74.845 248.045 74.905 ;
        RECT 258.765 75.045 259.085 75.105 ;
        RECT 260.695 75.090 260.835 75.245 ;
        RECT 261.065 75.185 261.385 75.245 ;
        RECT 260.160 75.045 260.450 75.090 ;
        RECT 258.765 74.905 260.450 75.045 ;
        RECT 258.765 74.845 259.085 74.905 ;
        RECT 260.160 74.860 260.450 74.905 ;
        RECT 260.625 74.860 260.915 75.090 ;
        RECT 261.525 74.845 261.845 75.105 ;
        RECT 262.075 75.045 262.215 75.585 ;
        RECT 262.445 75.585 263.685 75.725 ;
        RECT 262.445 75.525 262.765 75.585 ;
        RECT 263.365 75.525 263.685 75.585 ;
        RECT 281.880 75.725 282.170 75.770 ;
        RECT 285.000 75.725 285.290 75.770 ;
        RECT 286.890 75.725 287.180 75.770 ;
        RECT 281.880 75.585 287.180 75.725 ;
        RECT 281.880 75.540 282.170 75.585 ;
        RECT 285.000 75.540 285.290 75.585 ;
        RECT 286.890 75.540 287.180 75.585 ;
        RECT 295.530 75.725 295.820 75.770 ;
        RECT 297.420 75.725 297.710 75.770 ;
        RECT 300.540 75.725 300.830 75.770 ;
        RECT 295.530 75.585 300.830 75.725 ;
        RECT 295.530 75.540 295.820 75.585 ;
        RECT 297.420 75.540 297.710 75.585 ;
        RECT 300.540 75.540 300.830 75.585 ;
        RECT 276.245 75.185 276.565 75.445 ;
        RECT 277.180 75.385 277.470 75.430 ;
        RECT 283.145 75.385 283.465 75.445 ;
        RECT 277.180 75.245 283.465 75.385 ;
        RECT 277.180 75.200 277.470 75.245 ;
        RECT 283.145 75.185 283.465 75.245 ;
        RECT 287.760 75.385 288.050 75.430 ;
        RECT 290.505 75.385 290.825 75.445 ;
        RECT 293.280 75.385 293.570 75.430 ;
        RECT 287.760 75.245 293.570 75.385 ;
        RECT 287.760 75.200 288.050 75.245 ;
        RECT 290.505 75.185 290.825 75.245 ;
        RECT 293.280 75.200 293.570 75.245 ;
        RECT 298.325 75.385 298.645 75.445 ;
        RECT 298.325 75.245 302.235 75.385 ;
        RECT 298.325 75.185 298.645 75.245 ;
        RECT 262.690 75.045 262.980 75.090 ;
        RECT 264.285 75.045 264.605 75.105 ;
        RECT 262.075 74.905 268.655 75.045 ;
        RECT 262.690 74.860 262.980 74.905 ;
        RECT 264.285 74.845 264.605 74.905 ;
        RECT 212.305 74.750 212.625 74.765 ;
        RECT 208.740 74.705 209.330 74.750 ;
        RECT 211.980 74.705 212.630 74.750 ;
        RECT 208.740 74.565 212.630 74.705 ;
        RECT 208.740 74.520 209.030 74.565 ;
        RECT 211.980 74.520 212.630 74.565 ;
        RECT 214.620 74.705 214.910 74.750 ;
        RECT 216.905 74.705 217.225 74.765 ;
        RECT 214.620 74.565 217.225 74.705 ;
        RECT 214.620 74.520 214.910 74.565 ;
        RECT 212.305 74.505 212.625 74.520 ;
        RECT 216.905 74.505 217.225 74.565 ;
        RECT 219.205 74.505 219.525 74.765 ;
        RECT 241.285 74.705 241.605 74.765 ;
        RECT 243.585 74.705 243.905 74.765 ;
        RECT 241.285 74.565 243.905 74.705 ;
        RECT 241.285 74.505 241.605 74.565 ;
        RECT 243.585 74.505 243.905 74.565 ;
        RECT 257.845 74.705 258.165 74.765 ;
        RECT 262.000 74.705 262.290 74.750 ;
        RECT 267.965 74.705 268.285 74.765 ;
        RECT 257.845 74.565 268.285 74.705 ;
        RECT 268.515 74.705 268.655 74.905 ;
        RECT 275.785 74.845 276.105 75.105 ;
        RECT 277.165 74.705 277.485 74.765 ;
        RECT 268.515 74.565 277.485 74.705 ;
        RECT 257.845 74.505 258.165 74.565 ;
        RECT 262.000 74.520 262.290 74.565 ;
        RECT 267.965 74.505 268.285 74.565 ;
        RECT 277.165 74.505 277.485 74.565 ;
        RECT 277.640 74.705 277.930 74.750 ;
        RECT 278.085 74.705 278.405 74.765 ;
        RECT 280.800 74.750 281.090 75.065 ;
        RECT 281.880 75.045 282.170 75.090 ;
        RECT 285.460 75.045 285.750 75.090 ;
        RECT 287.295 75.045 287.585 75.090 ;
        RECT 281.880 74.905 287.585 75.045 ;
        RECT 281.880 74.860 282.170 74.905 ;
        RECT 285.460 74.860 285.750 74.905 ;
        RECT 287.295 74.860 287.585 74.905 ;
        RECT 288.205 75.045 288.525 75.105 ;
        RECT 289.585 75.045 289.905 75.105 ;
        RECT 288.205 74.905 289.905 75.045 ;
        RECT 288.205 74.845 288.525 74.905 ;
        RECT 289.585 74.845 289.905 74.905 ;
        RECT 294.645 74.845 294.965 75.105 ;
        RECT 295.125 75.045 295.415 75.090 ;
        RECT 296.960 75.045 297.250 75.090 ;
        RECT 300.540 75.045 300.830 75.090 ;
        RECT 295.125 74.905 300.830 75.045 ;
        RECT 295.125 74.860 295.415 74.905 ;
        RECT 296.960 74.860 297.250 74.905 ;
        RECT 300.540 74.860 300.830 74.905 ;
        RECT 284.065 74.750 284.385 74.765 ;
        RECT 277.640 74.565 278.405 74.705 ;
        RECT 277.640 74.520 277.930 74.565 ;
        RECT 278.085 74.505 278.405 74.565 ;
        RECT 280.500 74.705 281.090 74.750 ;
        RECT 283.740 74.705 284.390 74.750 ;
        RECT 280.500 74.565 285.675 74.705 ;
        RECT 280.500 74.520 280.790 74.565 ;
        RECT 283.740 74.520 284.390 74.565 ;
        RECT 284.065 74.505 284.385 74.520 ;
        RECT 285.535 74.425 285.675 74.565 ;
        RECT 286.365 74.505 286.685 74.765 ;
        RECT 294.185 74.705 294.505 74.765 ;
        RECT 301.620 74.750 301.910 75.065 ;
        RECT 302.095 74.750 302.235 75.245 ;
        RECT 307.065 75.185 307.385 75.445 ;
        RECT 302.925 75.045 303.245 75.105 ;
        RECT 306.160 75.045 306.450 75.090 ;
        RECT 302.925 74.905 306.450 75.045 ;
        RECT 302.925 74.845 303.245 74.905 ;
        RECT 306.160 74.860 306.450 74.905 ;
        RECT 296.040 74.705 296.330 74.750 ;
        RECT 294.185 74.565 296.330 74.705 ;
        RECT 294.185 74.505 294.505 74.565 ;
        RECT 296.040 74.520 296.330 74.565 ;
        RECT 298.320 74.705 298.970 74.750 ;
        RECT 301.620 74.705 302.235 74.750 ;
        RECT 302.465 74.705 302.785 74.765 ;
        RECT 306.620 74.705 306.910 74.750 ;
        RECT 298.320 74.565 302.785 74.705 ;
        RECT 298.320 74.520 298.970 74.565 ;
        RECT 301.920 74.520 302.210 74.565 ;
        RECT 302.465 74.505 302.785 74.565 ;
        RECT 303.015 74.565 306.910 74.705 ;
        RECT 215.065 74.365 215.385 74.425 ;
        RECT 207.335 74.225 215.385 74.365 ;
        RECT 192.525 74.165 192.845 74.225 ;
        RECT 201.740 74.180 202.030 74.225 ;
        RECT 215.065 74.165 215.385 74.225 ;
        RECT 218.285 74.165 218.605 74.425 ;
        RECT 218.760 74.365 219.050 74.410 ;
        RECT 219.665 74.365 219.985 74.425 ;
        RECT 259.225 74.365 259.545 74.425 ;
        RECT 261.065 74.365 261.385 74.425 ;
        RECT 218.760 74.225 261.385 74.365 ;
        RECT 218.760 74.180 219.050 74.225 ;
        RECT 219.665 74.165 219.985 74.225 ;
        RECT 259.225 74.165 259.545 74.225 ;
        RECT 261.065 74.165 261.385 74.225 ;
        RECT 263.380 74.365 263.670 74.410 ;
        RECT 266.585 74.365 266.905 74.425 ;
        RECT 263.380 74.225 266.905 74.365 ;
        RECT 263.380 74.180 263.670 74.225 ;
        RECT 266.585 74.165 266.905 74.225 ;
        RECT 279.005 74.165 279.325 74.425 ;
        RECT 285.445 74.165 285.765 74.425 ;
        RECT 289.585 74.365 289.905 74.425 ;
        RECT 303.015 74.365 303.155 74.565 ;
        RECT 306.620 74.520 306.910 74.565 ;
        RECT 289.585 74.225 303.155 74.365 ;
        RECT 289.585 74.165 289.905 74.225 ;
        RECT 162.095 73.545 311.135 74.025 ;
        RECT 173.205 73.345 173.525 73.405 ;
        RECT 188.845 73.345 189.165 73.405 ;
        RECT 192.065 73.345 192.385 73.405 ;
        RECT 170.075 73.205 189.165 73.345 ;
        RECT 170.075 72.710 170.215 73.205 ;
        RECT 173.205 73.145 173.525 73.205 ;
        RECT 188.845 73.145 189.165 73.205 ;
        RECT 189.395 73.205 192.385 73.345 ;
        RECT 173.660 73.005 174.310 73.050 ;
        RECT 177.260 73.005 177.550 73.050 ;
        RECT 173.660 72.865 177.550 73.005 ;
        RECT 173.660 72.820 174.310 72.865 ;
        RECT 176.960 72.820 177.550 72.865 ;
        RECT 186.545 73.005 186.865 73.065 ;
        RECT 189.395 73.005 189.535 73.205 ;
        RECT 192.065 73.145 192.385 73.205 ;
        RECT 194.365 73.345 194.685 73.405 ;
        RECT 196.680 73.345 196.970 73.390 ;
        RECT 194.365 73.205 196.970 73.345 ;
        RECT 194.365 73.145 194.685 73.205 ;
        RECT 196.680 73.160 196.970 73.205 ;
        RECT 198.980 73.345 199.270 73.390 ;
        RECT 200.345 73.345 200.665 73.405 ;
        RECT 202.185 73.345 202.505 73.405 ;
        RECT 243.125 73.345 243.445 73.405 ;
        RECT 270.725 73.345 271.045 73.405 ;
        RECT 198.980 73.205 200.665 73.345 ;
        RECT 198.980 73.160 199.270 73.205 ;
        RECT 200.345 73.145 200.665 73.205 ;
        RECT 200.895 73.205 202.505 73.345 ;
        RECT 186.545 72.865 189.535 73.005 ;
        RECT 189.780 73.005 190.070 73.050 ;
        RECT 190.225 73.005 190.545 73.065 ;
        RECT 191.605 73.005 191.925 73.065 ;
        RECT 198.520 73.005 198.810 73.050 ;
        RECT 200.895 73.005 201.035 73.205 ;
        RECT 202.185 73.145 202.505 73.205 ;
        RECT 205.035 73.205 241.055 73.345 ;
        RECT 205.035 73.065 205.175 73.205 ;
        RECT 204.025 73.005 204.345 73.065 ;
        RECT 189.780 72.865 191.925 73.005 ;
        RECT 176.960 72.725 177.250 72.820 ;
        RECT 186.545 72.805 186.865 72.865 ;
        RECT 189.780 72.820 190.070 72.865 ;
        RECT 190.225 72.805 190.545 72.865 ;
        RECT 191.605 72.805 191.925 72.865 ;
        RECT 192.155 72.865 201.035 73.005 ;
        RECT 201.815 72.865 204.345 73.005 ;
        RECT 170.000 72.480 170.290 72.710 ;
        RECT 170.465 72.665 170.755 72.710 ;
        RECT 172.300 72.665 172.590 72.710 ;
        RECT 175.880 72.665 176.170 72.710 ;
        RECT 170.465 72.525 176.170 72.665 ;
        RECT 170.465 72.480 170.755 72.525 ;
        RECT 172.300 72.480 172.590 72.525 ;
        RECT 175.880 72.480 176.170 72.525 ;
        RECT 176.885 72.505 177.250 72.725 ;
        RECT 182.865 72.665 183.185 72.725 ;
        RECT 185.180 72.665 185.470 72.710 ;
        RECT 192.155 72.665 192.295 72.865 ;
        RECT 198.520 72.820 198.810 72.865 ;
        RECT 182.865 72.525 185.470 72.665 ;
        RECT 176.885 72.465 177.205 72.505 ;
        RECT 182.865 72.465 183.185 72.525 ;
        RECT 185.180 72.480 185.470 72.525 ;
        RECT 185.715 72.525 192.295 72.665 ;
        RECT 171.380 72.325 171.670 72.370 ;
        RECT 174.125 72.325 174.445 72.385 ;
        RECT 171.380 72.185 174.445 72.325 ;
        RECT 171.380 72.140 171.670 72.185 ;
        RECT 174.125 72.125 174.445 72.185 ;
        RECT 176.425 72.325 176.745 72.385 ;
        RECT 178.740 72.325 179.030 72.370 ;
        RECT 176.425 72.185 179.030 72.325 ;
        RECT 176.425 72.125 176.745 72.185 ;
        RECT 178.740 72.140 179.030 72.185 ;
        RECT 181.025 72.325 181.345 72.385 ;
        RECT 185.715 72.325 185.855 72.525 ;
        RECT 193.445 72.465 193.765 72.725 ;
        RECT 201.815 72.710 201.955 72.865 ;
        RECT 204.025 72.805 204.345 72.865 ;
        RECT 204.945 72.805 205.265 73.065 ;
        RECT 210.465 73.005 210.785 73.065 ;
        RECT 219.205 73.005 219.525 73.065 ;
        RECT 221.965 73.050 222.285 73.065 ;
        RECT 210.465 72.865 216.215 73.005 ;
        RECT 210.465 72.805 210.785 72.865 ;
        RECT 195.835 72.525 201.495 72.665 ;
        RECT 181.025 72.185 185.855 72.325 ;
        RECT 187.925 72.325 188.245 72.385 ;
        RECT 195.835 72.325 195.975 72.525 ;
        RECT 187.925 72.185 195.975 72.325 ;
        RECT 181.025 72.125 181.345 72.185 ;
        RECT 187.925 72.125 188.245 72.185 ;
        RECT 199.900 72.140 200.190 72.370 ;
        RECT 170.870 71.985 171.160 72.030 ;
        RECT 172.760 71.985 173.050 72.030 ;
        RECT 175.880 71.985 176.170 72.030 ;
        RECT 170.870 71.845 176.170 71.985 ;
        RECT 199.975 71.985 200.115 72.140 ;
        RECT 200.805 72.125 201.125 72.385 ;
        RECT 201.355 72.325 201.495 72.525 ;
        RECT 201.740 72.480 202.030 72.710 ;
        RECT 203.580 72.665 203.870 72.710 ;
        RECT 208.165 72.665 208.485 72.725 ;
        RECT 203.580 72.525 208.485 72.665 ;
        RECT 203.580 72.480 203.870 72.525 ;
        RECT 203.655 72.325 203.795 72.480 ;
        RECT 208.165 72.465 208.485 72.525 ;
        RECT 211.400 72.480 211.690 72.710 ;
        RECT 211.860 72.665 212.150 72.710 ;
        RECT 215.065 72.665 215.385 72.725 ;
        RECT 216.075 72.710 216.215 72.865 ;
        RECT 217.915 72.865 219.525 73.005 ;
        RECT 211.860 72.525 215.385 72.665 ;
        RECT 211.860 72.480 212.150 72.525 ;
        RECT 201.355 72.185 203.795 72.325 ;
        RECT 204.025 72.325 204.345 72.385 ;
        RECT 210.925 72.325 211.245 72.385 ;
        RECT 211.475 72.325 211.615 72.480 ;
        RECT 215.065 72.465 215.385 72.525 ;
        RECT 215.540 72.480 215.830 72.710 ;
        RECT 216.000 72.480 216.290 72.710 ;
        RECT 216.460 72.480 216.750 72.710 ;
        RECT 204.025 72.185 211.615 72.325 ;
        RECT 212.780 72.325 213.070 72.370 ;
        RECT 213.225 72.325 213.545 72.385 ;
        RECT 212.780 72.185 213.545 72.325 ;
        RECT 204.025 72.125 204.345 72.185 ;
        RECT 210.925 72.125 211.245 72.185 ;
        RECT 212.780 72.140 213.070 72.185 ;
        RECT 203.120 71.985 203.410 72.030 ;
        RECT 203.565 71.985 203.885 72.045 ;
        RECT 199.975 71.845 203.885 71.985 ;
        RECT 170.870 71.800 171.160 71.845 ;
        RECT 172.760 71.800 173.050 71.845 ;
        RECT 175.880 71.800 176.170 71.845 ;
        RECT 203.120 71.800 203.410 71.845 ;
        RECT 203.565 71.785 203.885 71.845 ;
        RECT 204.485 71.985 204.805 72.045 ;
        RECT 212.855 71.985 212.995 72.140 ;
        RECT 213.225 72.125 213.545 72.185 ;
        RECT 214.145 72.125 214.465 72.385 ;
        RECT 214.605 72.325 214.925 72.385 ;
        RECT 215.615 72.325 215.755 72.480 ;
        RECT 214.605 72.185 215.755 72.325 ;
        RECT 214.605 72.125 214.925 72.185 ;
        RECT 204.485 71.845 212.995 71.985 ;
        RECT 204.485 71.785 204.805 71.845 ;
        RECT 171.825 71.645 172.145 71.705 ;
        RECT 177.345 71.645 177.665 71.705 ;
        RECT 204.025 71.645 204.345 71.705 ;
        RECT 171.825 71.505 204.345 71.645 ;
        RECT 171.825 71.445 172.145 71.505 ;
        RECT 177.345 71.445 177.665 71.505 ;
        RECT 204.025 71.445 204.345 71.505 ;
        RECT 208.625 71.645 208.945 71.705 ;
        RECT 209.560 71.645 209.850 71.690 ;
        RECT 208.625 71.505 209.850 71.645 ;
        RECT 208.625 71.445 208.945 71.505 ;
        RECT 209.560 71.460 209.850 71.505 ;
        RECT 213.225 71.645 213.545 71.705 ;
        RECT 216.535 71.645 216.675 72.480 ;
        RECT 217.365 72.465 217.685 72.725 ;
        RECT 217.915 72.710 218.055 72.865 ;
        RECT 219.205 72.805 219.525 72.865 ;
        RECT 221.500 73.005 222.285 73.050 ;
        RECT 225.100 73.005 225.390 73.050 ;
        RECT 221.500 72.865 225.390 73.005 ;
        RECT 221.500 72.820 222.285 72.865 ;
        RECT 221.965 72.805 222.285 72.820 ;
        RECT 224.800 72.820 225.390 72.865 ;
        RECT 227.485 73.005 227.805 73.065 ;
        RECT 227.485 72.865 231.855 73.005 ;
        RECT 217.840 72.480 218.130 72.710 ;
        RECT 218.305 72.665 218.595 72.710 ;
        RECT 220.140 72.665 220.430 72.710 ;
        RECT 223.720 72.665 224.010 72.710 ;
        RECT 218.305 72.525 224.010 72.665 ;
        RECT 218.305 72.480 218.595 72.525 ;
        RECT 220.140 72.480 220.430 72.525 ;
        RECT 223.720 72.480 224.010 72.525 ;
        RECT 224.800 72.505 225.090 72.820 ;
        RECT 227.485 72.805 227.805 72.865 ;
        RECT 229.785 72.465 230.105 72.725 ;
        RECT 230.705 72.465 231.025 72.725 ;
        RECT 231.165 72.465 231.485 72.725 ;
        RECT 231.715 72.710 231.855 72.865 ;
        RECT 240.915 72.725 241.055 73.205 ;
        RECT 243.125 73.205 271.045 73.345 ;
        RECT 243.125 73.145 243.445 73.205 ;
        RECT 270.725 73.145 271.045 73.205 ;
        RECT 283.605 73.345 283.925 73.405 ;
        RECT 287.300 73.345 287.590 73.390 ;
        RECT 283.605 73.205 287.590 73.345 ;
        RECT 283.605 73.145 283.925 73.205 ;
        RECT 287.300 73.160 287.590 73.205 ;
        RECT 302.925 73.345 303.245 73.405 ;
        RECT 304.320 73.345 304.610 73.390 ;
        RECT 302.925 73.205 304.610 73.345 ;
        RECT 302.925 73.145 303.245 73.205 ;
        RECT 304.320 73.160 304.610 73.205 ;
        RECT 241.745 72.805 242.065 73.065 ;
        RECT 244.980 73.005 245.270 73.050 ;
        RECT 250.025 73.005 250.345 73.065 ;
        RECT 259.225 73.005 259.545 73.065 ;
        RECT 261.540 73.005 261.830 73.050 ;
        RECT 263.365 73.005 263.685 73.065 ;
        RECT 244.980 72.865 250.345 73.005 ;
        RECT 244.980 72.820 245.270 72.865 ;
        RECT 250.025 72.805 250.345 72.865 ;
        RECT 255.865 72.865 259.915 73.005 ;
        RECT 231.640 72.480 231.930 72.710 ;
        RECT 234.385 72.665 234.705 72.725 ;
        RECT 239.920 72.665 240.210 72.710 ;
        RECT 234.385 72.525 240.210 72.665 ;
        RECT 234.385 72.465 234.705 72.525 ;
        RECT 239.920 72.480 240.210 72.525 ;
        RECT 240.385 72.480 240.675 72.710 ;
        RECT 240.825 72.665 241.145 72.725 ;
        RECT 241.300 72.665 241.590 72.710 ;
        RECT 240.825 72.525 241.590 72.665 ;
        RECT 219.205 72.125 219.525 72.385 ;
        RECT 225.185 72.325 225.505 72.385 ;
        RECT 226.580 72.325 226.870 72.370 ;
        RECT 240.460 72.325 240.600 72.480 ;
        RECT 240.825 72.465 241.145 72.525 ;
        RECT 241.300 72.480 241.590 72.525 ;
        RECT 242.450 72.480 242.740 72.710 ;
        RECT 243.585 72.665 243.905 72.725 ;
        RECT 245.885 72.710 246.205 72.725 ;
        RECT 244.290 72.665 244.580 72.710 ;
        RECT 243.585 72.525 244.580 72.665 ;
        RECT 225.185 72.185 240.600 72.325 ;
        RECT 242.525 72.325 242.665 72.480 ;
        RECT 243.585 72.465 243.905 72.525 ;
        RECT 244.290 72.480 244.580 72.525 ;
        RECT 245.440 72.480 245.730 72.710 ;
        RECT 245.885 72.480 246.370 72.710 ;
        RECT 246.805 72.665 247.125 72.725 ;
        RECT 255.865 72.665 256.005 72.865 ;
        RECT 259.225 72.805 259.545 72.865 ;
        RECT 246.805 72.525 256.005 72.665 ;
        RECT 245.515 72.325 245.655 72.480 ;
        RECT 245.885 72.465 246.205 72.480 ;
        RECT 246.805 72.465 247.125 72.525 ;
        RECT 256.465 72.465 256.785 72.725 ;
        RECT 257.400 72.480 257.690 72.710 ;
        RECT 252.785 72.325 253.105 72.385 ;
        RECT 242.525 72.185 244.270 72.325 ;
        RECT 245.515 72.185 253.105 72.325 ;
        RECT 225.185 72.125 225.505 72.185 ;
        RECT 226.580 72.140 226.870 72.185 ;
        RECT 218.710 71.985 219.000 72.030 ;
        RECT 220.600 71.985 220.890 72.030 ;
        RECT 223.720 71.985 224.010 72.030 ;
        RECT 218.710 71.845 224.010 71.985 ;
        RECT 218.710 71.800 219.000 71.845 ;
        RECT 220.600 71.800 220.890 71.845 ;
        RECT 223.720 71.800 224.010 71.845 ;
        RECT 230.705 71.985 231.025 72.045 ;
        RECT 232.085 71.985 232.405 72.045 ;
        RECT 230.705 71.845 232.405 71.985 ;
        RECT 230.705 71.785 231.025 71.845 ;
        RECT 232.085 71.785 232.405 71.845 ;
        RECT 241.745 71.985 242.065 72.045 ;
        RECT 243.600 71.985 243.890 72.030 ;
        RECT 241.745 71.845 243.890 71.985 ;
        RECT 244.130 71.985 244.270 72.185 ;
        RECT 252.785 72.125 253.105 72.185 ;
        RECT 253.245 72.325 253.565 72.385 ;
        RECT 257.475 72.325 257.615 72.480 ;
        RECT 257.845 72.465 258.165 72.725 ;
        RECT 258.305 72.465 258.625 72.725 ;
        RECT 259.775 72.710 259.915 72.865 ;
        RECT 261.540 72.865 263.685 73.005 ;
        RECT 261.540 72.820 261.830 72.865 ;
        RECT 263.365 72.805 263.685 72.865 ;
        RECT 265.665 73.005 265.985 73.065 ;
        RECT 267.520 73.005 267.810 73.050 ;
        RECT 272.105 73.005 272.425 73.065 ;
        RECT 265.665 72.865 272.425 73.005 ;
        RECT 265.665 72.805 265.985 72.865 ;
        RECT 267.520 72.820 267.810 72.865 ;
        RECT 272.105 72.805 272.425 72.865 ;
        RECT 279.925 72.805 280.245 73.065 ;
        RECT 282.220 73.005 282.870 73.050 ;
        RECT 285.820 73.005 286.110 73.050 ;
        RECT 282.220 72.865 286.110 73.005 ;
        RECT 282.220 72.820 282.870 72.865 ;
        RECT 285.520 72.820 286.110 72.865 ;
        RECT 285.520 72.725 285.810 72.820 ;
        RECT 290.505 72.805 290.825 73.065 ;
        RECT 298.325 73.050 298.645 73.065 ;
        RECT 294.760 73.005 295.050 73.050 ;
        RECT 298.000 73.005 298.650 73.050 ;
        RECT 299.245 73.005 299.565 73.065 ;
        RECT 294.760 72.865 299.565 73.005 ;
        RECT 294.760 72.820 295.350 72.865 ;
        RECT 298.000 72.820 298.650 72.865 ;
        RECT 260.605 72.710 260.925 72.725 ;
        RECT 259.700 72.480 259.990 72.710 ;
        RECT 260.440 72.480 260.925 72.710 ;
        RECT 261.080 72.665 261.370 72.710 ;
        RECT 262.220 72.665 262.510 72.710 ;
        RECT 264.285 72.665 264.605 72.725 ;
        RECT 261.080 72.525 261.755 72.665 ;
        RECT 261.080 72.480 261.370 72.525 ;
        RECT 260.605 72.465 260.925 72.480 ;
        RECT 253.245 72.185 257.615 72.325 ;
        RECT 253.245 72.125 253.565 72.185 ;
        RECT 249.105 71.985 249.425 72.045 ;
        RECT 254.625 71.985 254.945 72.045 ;
        RECT 258.305 71.985 258.625 72.045 ;
        RECT 261.615 71.985 261.755 72.525 ;
        RECT 262.220 72.525 264.605 72.665 ;
        RECT 262.220 72.480 262.510 72.525 ;
        RECT 264.285 72.465 264.605 72.525 ;
        RECT 265.205 72.665 265.525 72.725 ;
        RECT 266.600 72.665 266.890 72.710 ;
        RECT 265.205 72.525 266.890 72.665 ;
        RECT 265.205 72.465 265.525 72.525 ;
        RECT 266.600 72.480 266.890 72.525 ;
        RECT 267.060 72.665 267.350 72.710 ;
        RECT 267.965 72.665 268.285 72.725 ;
        RECT 267.060 72.525 268.285 72.665 ;
        RECT 267.060 72.480 267.350 72.525 ;
        RECT 267.965 72.465 268.285 72.525 ;
        RECT 268.440 72.665 268.730 72.710 ;
        RECT 268.885 72.665 269.205 72.725 ;
        RECT 268.440 72.525 269.205 72.665 ;
        RECT 268.440 72.480 268.730 72.525 ;
        RECT 268.885 72.465 269.205 72.525 ;
        RECT 277.180 72.665 277.470 72.710 ;
        RECT 278.085 72.665 278.405 72.725 ;
        RECT 277.180 72.525 278.405 72.665 ;
        RECT 277.180 72.480 277.470 72.525 ;
        RECT 278.085 72.465 278.405 72.525 ;
        RECT 279.025 72.665 279.315 72.710 ;
        RECT 280.860 72.665 281.150 72.710 ;
        RECT 284.440 72.665 284.730 72.710 ;
        RECT 279.025 72.525 284.730 72.665 ;
        RECT 279.025 72.480 279.315 72.525 ;
        RECT 280.860 72.480 281.150 72.525 ;
        RECT 284.440 72.480 284.730 72.525 ;
        RECT 285.445 72.665 285.810 72.725 ;
        RECT 286.825 72.665 287.145 72.725 ;
        RECT 285.445 72.525 287.145 72.665 ;
        RECT 285.445 72.505 285.810 72.525 ;
        RECT 285.445 72.465 285.765 72.505 ;
        RECT 286.825 72.465 287.145 72.525 ;
        RECT 295.060 72.505 295.350 72.820 ;
        RECT 298.325 72.805 298.645 72.820 ;
        RECT 299.245 72.805 299.565 72.865 ;
        RECT 300.640 73.005 300.930 73.050 ;
        RECT 300.640 72.865 302.235 73.005 ;
        RECT 300.640 72.820 300.930 72.865 ;
        RECT 296.140 72.665 296.430 72.710 ;
        RECT 299.720 72.665 300.010 72.710 ;
        RECT 301.555 72.665 301.845 72.710 ;
        RECT 296.140 72.525 301.845 72.665 ;
        RECT 302.095 72.665 302.235 72.865 ;
        RECT 307.065 72.665 307.385 72.725 ;
        RECT 302.095 72.525 302.695 72.665 ;
        RECT 296.140 72.480 296.430 72.525 ;
        RECT 299.720 72.480 300.010 72.525 ;
        RECT 301.555 72.480 301.845 72.525 ;
        RECT 275.800 72.325 276.090 72.370 ;
        RECT 276.245 72.325 276.565 72.385 ;
        RECT 244.130 71.845 258.625 71.985 ;
        RECT 241.745 71.785 242.065 71.845 ;
        RECT 243.600 71.800 243.890 71.845 ;
        RECT 249.105 71.785 249.425 71.845 ;
        RECT 254.625 71.785 254.945 71.845 ;
        RECT 258.305 71.785 258.625 71.845 ;
        RECT 258.855 71.845 261.755 71.985 ;
        RECT 262.560 72.185 268.655 72.325 ;
        RECT 213.225 71.505 216.675 71.645 ;
        RECT 213.225 71.445 213.545 71.505 ;
        RECT 232.545 71.445 232.865 71.705 ;
        RECT 241.285 71.645 241.605 71.705 ;
        RECT 243.140 71.645 243.430 71.690 ;
        RECT 241.285 71.505 243.430 71.645 ;
        RECT 241.285 71.445 241.605 71.505 ;
        RECT 243.140 71.460 243.430 71.505 ;
        RECT 253.705 71.645 254.025 71.705 ;
        RECT 258.855 71.645 258.995 71.845 ;
        RECT 253.705 71.505 258.995 71.645 ;
        RECT 259.240 71.645 259.530 71.690 ;
        RECT 262.560 71.645 262.700 72.185 ;
        RECT 268.515 72.045 268.655 72.185 ;
        RECT 275.800 72.185 276.565 72.325 ;
        RECT 275.800 72.140 276.090 72.185 ;
        RECT 276.245 72.125 276.565 72.185 ;
        RECT 278.545 72.125 278.865 72.385 ;
        RECT 294.645 72.325 294.965 72.385 ;
        RECT 302.020 72.325 302.310 72.370 ;
        RECT 294.645 72.185 302.310 72.325 ;
        RECT 294.645 72.125 294.965 72.185 ;
        RECT 302.020 72.140 302.310 72.185 ;
        RECT 262.920 71.985 263.210 72.030 ;
        RECT 267.505 71.985 267.825 72.045 ;
        RECT 262.920 71.845 267.825 71.985 ;
        RECT 262.920 71.800 263.210 71.845 ;
        RECT 267.505 71.785 267.825 71.845 ;
        RECT 268.425 71.785 268.745 72.045 ;
        RECT 302.555 72.030 302.695 72.525 ;
        RECT 304.395 72.525 307.385 72.665 ;
        RECT 303.385 72.325 303.705 72.385 ;
        RECT 304.395 72.325 304.535 72.525 ;
        RECT 305.315 72.370 305.455 72.525 ;
        RECT 307.065 72.465 307.385 72.525 ;
        RECT 307.525 72.665 307.845 72.725 ;
        RECT 308.000 72.665 308.290 72.710 ;
        RECT 307.525 72.525 308.290 72.665 ;
        RECT 307.525 72.465 307.845 72.525 ;
        RECT 308.000 72.480 308.290 72.525 ;
        RECT 303.385 72.185 304.535 72.325 ;
        RECT 303.385 72.125 303.705 72.185 ;
        RECT 304.780 72.140 305.070 72.370 ;
        RECT 305.240 72.140 305.530 72.370 ;
        RECT 279.430 71.985 279.720 72.030 ;
        RECT 281.320 71.985 281.610 72.030 ;
        RECT 284.440 71.985 284.730 72.030 ;
        RECT 279.430 71.845 284.730 71.985 ;
        RECT 279.430 71.800 279.720 71.845 ;
        RECT 281.320 71.800 281.610 71.845 ;
        RECT 284.440 71.800 284.730 71.845 ;
        RECT 296.140 71.985 296.430 72.030 ;
        RECT 299.260 71.985 299.550 72.030 ;
        RECT 301.150 71.985 301.440 72.030 ;
        RECT 296.140 71.845 301.440 71.985 ;
        RECT 296.140 71.800 296.430 71.845 ;
        RECT 299.260 71.800 299.550 71.845 ;
        RECT 301.150 71.800 301.440 71.845 ;
        RECT 302.480 71.800 302.770 72.030 ;
        RECT 259.240 71.505 262.700 71.645 ;
        RECT 253.705 71.445 254.025 71.505 ;
        RECT 259.240 71.460 259.530 71.505 ;
        RECT 265.665 71.445 265.985 71.705 ;
        RECT 272.105 71.645 272.425 71.705 ;
        RECT 276.260 71.645 276.550 71.690 ;
        RECT 272.105 71.505 276.550 71.645 ;
        RECT 272.105 71.445 272.425 71.505 ;
        RECT 276.260 71.460 276.550 71.505 ;
        RECT 278.100 71.645 278.390 71.690 ;
        RECT 290.965 71.645 291.285 71.705 ;
        RECT 278.100 71.505 291.285 71.645 ;
        RECT 278.100 71.460 278.390 71.505 ;
        RECT 290.965 71.445 291.285 71.505 ;
        RECT 293.265 71.445 293.585 71.705 ;
        RECT 295.565 71.645 295.885 71.705 ;
        RECT 304.855 71.645 304.995 72.140 ;
        RECT 295.565 71.505 304.995 71.645 ;
        RECT 305.225 71.645 305.545 71.705 ;
        RECT 307.080 71.645 307.370 71.690 ;
        RECT 305.225 71.505 307.370 71.645 ;
        RECT 295.565 71.445 295.885 71.505 ;
        RECT 305.225 71.445 305.545 71.505 ;
        RECT 307.080 71.460 307.370 71.505 ;
        RECT 162.095 70.825 311.135 71.305 ;
        RECT 164.925 70.625 165.245 70.685 ;
        RECT 187.005 70.625 187.325 70.685 ;
        RECT 164.925 70.485 187.325 70.625 ;
        RECT 164.925 70.425 165.245 70.485 ;
        RECT 164.465 70.285 164.785 70.345 ;
        RECT 164.465 70.145 173.895 70.285 ;
        RECT 164.465 70.085 164.785 70.145 ;
        RECT 166.765 69.945 167.085 70.005 ;
        RECT 172.285 69.945 172.605 70.005 ;
        RECT 173.220 69.945 173.510 69.990 ;
        RECT 166.765 69.805 173.510 69.945 ;
        RECT 166.765 69.745 167.085 69.805 ;
        RECT 172.285 69.745 172.605 69.805 ;
        RECT 173.220 69.760 173.510 69.805 ;
        RECT 173.755 69.605 173.895 70.145 ;
        RECT 174.140 69.945 174.430 69.990 ;
        RECT 178.740 69.945 179.030 69.990 ;
        RECT 179.645 69.945 179.965 70.005 ;
        RECT 174.140 69.805 179.965 69.945 ;
        RECT 174.140 69.760 174.430 69.805 ;
        RECT 178.740 69.760 179.030 69.805 ;
        RECT 179.645 69.745 179.965 69.805 ;
        RECT 177.805 69.605 178.125 69.665 ;
        RECT 173.755 69.465 178.125 69.605 ;
        RECT 177.805 69.405 178.125 69.465 ;
        RECT 183.785 69.405 184.105 69.665 ;
        RECT 184.335 69.605 184.475 70.485 ;
        RECT 187.005 70.425 187.325 70.485 ;
        RECT 187.465 70.625 187.785 70.685 ;
        RECT 187.940 70.625 188.230 70.670 ;
        RECT 187.465 70.485 188.230 70.625 ;
        RECT 187.465 70.425 187.785 70.485 ;
        RECT 187.940 70.440 188.230 70.485 ;
        RECT 188.385 70.425 188.705 70.685 ;
        RECT 190.225 70.625 190.545 70.685 ;
        RECT 209.545 70.625 209.865 70.685 ;
        RECT 214.605 70.625 214.925 70.685 ;
        RECT 190.225 70.485 214.925 70.625 ;
        RECT 190.225 70.425 190.545 70.485 ;
        RECT 209.545 70.425 209.865 70.485 ;
        RECT 214.605 70.425 214.925 70.485 ;
        RECT 215.525 70.625 215.845 70.685 ;
        RECT 216.000 70.625 216.290 70.670 ;
        RECT 217.825 70.625 218.145 70.685 ;
        RECT 215.525 70.485 216.290 70.625 ;
        RECT 215.525 70.425 215.845 70.485 ;
        RECT 216.000 70.440 216.290 70.485 ;
        RECT 216.995 70.485 218.145 70.625 ;
        RECT 185.180 70.285 185.470 70.330 ;
        RECT 185.625 70.285 185.945 70.345 ;
        RECT 192.065 70.285 192.385 70.345 ;
        RECT 185.180 70.145 185.945 70.285 ;
        RECT 185.180 70.100 185.470 70.145 ;
        RECT 185.625 70.085 185.945 70.145 ;
        RECT 191.235 70.145 192.385 70.285 ;
        RECT 184.720 69.945 185.010 69.990 ;
        RECT 186.560 69.945 186.850 69.990 ;
        RECT 184.720 69.805 190.455 69.945 ;
        RECT 184.720 69.760 185.010 69.805 ;
        RECT 186.560 69.760 186.850 69.805 ;
        RECT 185.165 69.650 185.485 69.665 ;
        RECT 185.150 69.605 185.485 69.650 ;
        RECT 184.335 69.465 185.485 69.605 ;
        RECT 185.150 69.420 185.485 69.465 ;
        RECT 185.165 69.405 185.485 69.420 ;
        RECT 186.085 69.405 186.405 69.665 ;
        RECT 187.005 69.405 187.325 69.665 ;
        RECT 190.315 69.605 190.455 69.805 ;
        RECT 190.685 69.745 191.005 70.005 ;
        RECT 191.235 69.990 191.375 70.145 ;
        RECT 192.065 70.085 192.385 70.145 ;
        RECT 208.130 70.285 208.420 70.330 ;
        RECT 210.020 70.285 210.310 70.330 ;
        RECT 213.140 70.285 213.430 70.330 ;
        RECT 208.130 70.145 213.430 70.285 ;
        RECT 208.130 70.100 208.420 70.145 ;
        RECT 210.020 70.100 210.310 70.145 ;
        RECT 213.140 70.100 213.430 70.145 ;
        RECT 191.160 69.760 191.450 69.990 ;
        RECT 207.260 69.945 207.550 69.990 ;
        RECT 211.845 69.945 212.165 70.005 ;
        RECT 216.995 69.990 217.135 70.485 ;
        RECT 217.825 70.425 218.145 70.485 ;
        RECT 219.205 70.625 219.525 70.685 ;
        RECT 220.140 70.625 220.430 70.670 ;
        RECT 260.145 70.625 260.465 70.685 ;
        RECT 219.205 70.485 220.430 70.625 ;
        RECT 219.205 70.425 219.525 70.485 ;
        RECT 220.140 70.440 220.430 70.485 ;
        RECT 221.365 70.485 260.465 70.625 ;
        RECT 217.365 70.285 217.685 70.345 ;
        RECT 221.365 70.285 221.505 70.485 ;
        RECT 260.145 70.425 260.465 70.485 ;
        RECT 260.620 70.625 260.910 70.670 ;
        RECT 260.620 70.485 265.435 70.625 ;
        RECT 260.620 70.440 260.910 70.485 ;
        RECT 217.365 70.145 221.505 70.285 ;
        RECT 227.025 70.285 227.345 70.345 ;
        RECT 232.085 70.285 232.405 70.345 ;
        RECT 263.840 70.285 264.130 70.330 ;
        RECT 227.025 70.145 232.405 70.285 ;
        RECT 217.365 70.085 217.685 70.145 ;
        RECT 227.025 70.085 227.345 70.145 ;
        RECT 232.085 70.085 232.405 70.145 ;
        RECT 232.635 70.145 258.995 70.285 ;
        RECT 207.260 69.805 212.165 69.945 ;
        RECT 207.260 69.760 207.550 69.805 ;
        RECT 211.845 69.745 212.165 69.805 ;
        RECT 216.920 69.760 217.210 69.990 ;
        RECT 231.625 69.945 231.945 70.005 ;
        RECT 217.455 69.805 231.945 69.945 ;
        RECT 217.455 69.665 217.595 69.805 ;
        RECT 231.625 69.745 231.945 69.805 ;
        RECT 193.460 69.605 193.750 69.650 ;
        RECT 194.365 69.605 194.685 69.665 ;
        RECT 190.315 69.465 194.685 69.605 ;
        RECT 193.460 69.420 193.750 69.465 ;
        RECT 194.365 69.405 194.685 69.465 ;
        RECT 195.300 69.420 195.590 69.650 ;
        RECT 197.600 69.605 197.890 69.650 ;
        RECT 200.345 69.605 200.665 69.665 ;
        RECT 197.600 69.465 200.665 69.605 ;
        RECT 197.600 69.420 197.890 69.465 ;
        RECT 181.025 69.265 181.345 69.325 ;
        RECT 180.195 69.125 181.345 69.265 ;
        RECT 187.095 69.265 187.235 69.405 ;
        RECT 195.375 69.265 195.515 69.420 ;
        RECT 200.345 69.405 200.665 69.465 ;
        RECT 207.725 69.605 208.015 69.650 ;
        RECT 209.560 69.605 209.850 69.650 ;
        RECT 213.140 69.605 213.430 69.650 ;
        RECT 207.725 69.465 213.430 69.605 ;
        RECT 207.725 69.420 208.015 69.465 ;
        RECT 209.560 69.420 209.850 69.465 ;
        RECT 213.140 69.420 213.430 69.465 ;
        RECT 195.745 69.265 196.065 69.325 ;
        RECT 187.095 69.125 196.065 69.265 ;
        RECT 168.605 68.925 168.925 68.985 ;
        RECT 170.920 68.925 171.210 68.970 ;
        RECT 168.605 68.785 171.210 68.925 ;
        RECT 168.605 68.725 168.925 68.785 ;
        RECT 170.920 68.740 171.210 68.785 ;
        RECT 171.825 68.925 172.145 68.985 ;
        RECT 172.760 68.925 173.050 68.970 ;
        RECT 171.825 68.785 173.050 68.925 ;
        RECT 171.825 68.725 172.145 68.785 ;
        RECT 172.760 68.740 173.050 68.785 ;
        RECT 175.505 68.725 175.825 68.985 ;
        RECT 176.425 68.925 176.745 68.985 ;
        RECT 177.360 68.925 177.650 68.970 ;
        RECT 180.195 68.925 180.335 69.125 ;
        RECT 181.025 69.065 181.345 69.125 ;
        RECT 195.745 69.065 196.065 69.125 ;
        RECT 200.805 69.265 201.125 69.325 ;
        RECT 200.805 69.125 207.705 69.265 ;
        RECT 200.805 69.065 201.125 69.125 ;
        RECT 176.425 68.785 180.335 68.925 ;
        RECT 190.225 68.925 190.545 68.985 ;
        RECT 193.905 68.925 194.225 68.985 ;
        RECT 190.225 68.785 194.225 68.925 ;
        RECT 176.425 68.725 176.745 68.785 ;
        RECT 177.360 68.740 177.650 68.785 ;
        RECT 190.225 68.725 190.545 68.785 ;
        RECT 193.905 68.725 194.225 68.785 ;
        RECT 197.140 68.925 197.430 68.970 ;
        RECT 204.945 68.925 205.265 68.985 ;
        RECT 197.140 68.785 205.265 68.925 ;
        RECT 207.565 68.925 207.705 69.125 ;
        RECT 208.625 69.065 208.945 69.325 ;
        RECT 210.920 69.265 211.570 69.310 ;
        RECT 212.305 69.265 212.625 69.325 ;
        RECT 214.220 69.310 214.510 69.625 ;
        RECT 217.365 69.405 217.685 69.665 ;
        RECT 217.840 69.605 218.130 69.650 ;
        RECT 225.185 69.605 225.505 69.665 ;
        RECT 217.840 69.465 225.505 69.605 ;
        RECT 217.840 69.420 218.130 69.465 ;
        RECT 225.185 69.405 225.505 69.465 ;
        RECT 230.705 69.605 231.025 69.665 ;
        RECT 232.635 69.605 232.775 70.145 ;
        RECT 234.385 69.745 234.705 70.005 ;
        RECT 244.505 69.945 244.825 70.005 ;
        RECT 256.005 69.945 256.325 70.005 ;
        RECT 258.855 69.945 258.995 70.145 ;
        RECT 263.840 70.145 264.975 70.285 ;
        RECT 263.840 70.100 264.130 70.145 ;
        RECT 261.525 69.945 261.845 70.005 ;
        RECT 244.505 69.805 247.495 69.945 ;
        RECT 244.505 69.745 244.825 69.805 ;
        RECT 230.705 69.465 232.775 69.605 ;
        RECT 235.780 69.605 236.070 69.650 ;
        RECT 236.225 69.605 236.545 69.665 ;
        RECT 235.780 69.465 236.545 69.605 ;
        RECT 230.705 69.405 231.025 69.465 ;
        RECT 235.780 69.420 236.070 69.465 ;
        RECT 236.225 69.405 236.545 69.465 ;
        RECT 238.985 69.605 239.305 69.665 ;
        RECT 240.365 69.605 240.685 69.665 ;
        RECT 238.985 69.465 240.685 69.605 ;
        RECT 238.985 69.405 239.305 69.465 ;
        RECT 240.365 69.405 240.685 69.465 ;
        RECT 245.425 69.605 245.745 69.665 ;
        RECT 246.335 69.650 247.035 69.655 ;
        RECT 247.355 69.650 247.495 69.805 ;
        RECT 256.005 69.805 258.075 69.945 ;
        RECT 256.005 69.745 256.325 69.805 ;
        RECT 246.335 69.605 247.110 69.650 ;
        RECT 245.425 69.515 247.110 69.605 ;
        RECT 245.425 69.465 246.475 69.515 ;
        RECT 245.425 69.405 245.745 69.465 ;
        RECT 246.820 69.420 247.110 69.515 ;
        RECT 247.285 69.420 247.575 69.650 ;
        RECT 248.185 69.405 248.505 69.665 ;
        RECT 248.645 69.405 248.965 69.665 ;
        RECT 249.105 69.650 249.425 69.665 ;
        RECT 249.105 69.605 249.435 69.650 ;
        RECT 249.105 69.465 249.620 69.605 ;
        RECT 249.105 69.420 249.435 69.465 ;
        RECT 249.105 69.405 249.425 69.420 ;
        RECT 257.385 69.405 257.705 69.665 ;
        RECT 257.935 69.650 258.075 69.805 ;
        RECT 258.855 69.805 261.845 69.945 ;
        RECT 258.855 69.650 258.995 69.805 ;
        RECT 261.525 69.745 261.845 69.805 ;
        RECT 261.985 69.745 262.305 70.005 ;
        RECT 264.285 69.945 264.605 70.005 ;
        RECT 264.835 69.990 264.975 70.145 ;
        RECT 262.995 69.805 264.605 69.945 ;
        RECT 257.865 69.420 258.155 69.650 ;
        RECT 258.780 69.420 259.070 69.650 ;
        RECT 259.225 69.405 259.545 69.665 ;
        RECT 259.685 69.650 260.005 69.665 ;
        RECT 259.685 69.605 260.015 69.650 ;
        RECT 259.685 69.465 260.200 69.605 ;
        RECT 259.685 69.420 260.015 69.465 ;
        RECT 259.685 69.405 260.005 69.420 ;
        RECT 261.065 69.405 261.385 69.665 ;
        RECT 262.075 69.605 262.215 69.745 ;
        RECT 262.995 69.650 263.135 69.805 ;
        RECT 264.285 69.745 264.605 69.805 ;
        RECT 264.760 69.760 265.050 69.990 ;
        RECT 265.295 69.945 265.435 70.485 ;
        RECT 265.665 70.425 265.985 70.685 ;
        RECT 267.505 70.425 267.825 70.685 ;
        RECT 267.965 70.625 268.285 70.685 ;
        RECT 285.905 70.625 286.225 70.685 ;
        RECT 267.965 70.485 286.225 70.625 ;
        RECT 267.965 70.425 268.285 70.485 ;
        RECT 285.905 70.425 286.225 70.485 ;
        RECT 286.365 70.625 286.685 70.685 ;
        RECT 288.220 70.625 288.510 70.670 ;
        RECT 286.365 70.485 288.510 70.625 ;
        RECT 286.365 70.425 286.685 70.485 ;
        RECT 288.220 70.440 288.510 70.485 ;
        RECT 304.320 70.625 304.610 70.670 ;
        RECT 304.765 70.625 305.085 70.685 ;
        RECT 304.320 70.485 305.085 70.625 ;
        RECT 304.320 70.440 304.610 70.485 ;
        RECT 304.765 70.425 305.085 70.485 ;
        RECT 279.430 70.285 279.720 70.330 ;
        RECT 281.320 70.285 281.610 70.330 ;
        RECT 284.440 70.285 284.730 70.330 ;
        RECT 295.530 70.285 295.820 70.330 ;
        RECT 297.420 70.285 297.710 70.330 ;
        RECT 300.540 70.285 300.830 70.330 ;
        RECT 279.430 70.145 284.730 70.285 ;
        RECT 279.430 70.100 279.720 70.145 ;
        RECT 281.320 70.100 281.610 70.145 ;
        RECT 284.440 70.100 284.730 70.145 ;
        RECT 286.455 70.145 291.195 70.285 ;
        RECT 267.980 69.945 268.270 69.990 ;
        RECT 265.295 69.805 268.270 69.945 ;
        RECT 267.980 69.760 268.270 69.805 ;
        RECT 272.105 69.745 272.425 70.005 ;
        RECT 283.145 69.945 283.465 70.005 ;
        RECT 286.455 69.945 286.595 70.145 ;
        RECT 283.145 69.805 286.595 69.945 ;
        RECT 287.745 69.945 288.065 70.005 ;
        RECT 291.055 69.990 291.195 70.145 ;
        RECT 295.530 70.145 300.830 70.285 ;
        RECT 295.530 70.100 295.820 70.145 ;
        RECT 297.420 70.100 297.710 70.145 ;
        RECT 300.540 70.100 300.830 70.145 ;
        RECT 290.520 69.945 290.810 69.990 ;
        RECT 287.745 69.805 290.810 69.945 ;
        RECT 283.145 69.745 283.465 69.805 ;
        RECT 287.745 69.745 288.065 69.805 ;
        RECT 290.520 69.760 290.810 69.805 ;
        RECT 290.980 69.760 291.270 69.990 ;
        RECT 307.065 69.745 307.385 70.005 ;
        RECT 262.460 69.605 262.750 69.650 ;
        RECT 262.075 69.465 262.750 69.605 ;
        RECT 262.460 69.420 262.750 69.465 ;
        RECT 262.920 69.420 263.210 69.650 ;
        RECT 263.825 69.605 264.145 69.665 ;
        RECT 265.680 69.605 265.970 69.650 ;
        RECT 266.585 69.605 266.905 69.665 ;
        RECT 263.825 69.465 265.970 69.605 ;
        RECT 214.220 69.265 214.810 69.310 ;
        RECT 210.920 69.125 214.810 69.265 ;
        RECT 210.920 69.080 211.570 69.125 ;
        RECT 212.305 69.065 212.625 69.125 ;
        RECT 214.520 69.080 214.810 69.125 ;
        RECT 237.160 69.265 237.450 69.310 ;
        RECT 244.505 69.265 244.825 69.325 ;
        RECT 237.160 69.125 244.825 69.265 ;
        RECT 237.160 69.080 237.450 69.125 ;
        RECT 244.505 69.065 244.825 69.125 ;
        RECT 246.345 69.065 246.665 69.325 ;
        RECT 253.705 69.265 254.025 69.325 ;
        RECT 253.705 69.125 261.755 69.265 ;
        RECT 253.705 69.065 254.025 69.125 ;
        RECT 217.365 68.925 217.685 68.985 ;
        RECT 207.565 68.785 217.685 68.925 ;
        RECT 197.140 68.740 197.430 68.785 ;
        RECT 204.945 68.725 205.265 68.785 ;
        RECT 217.365 68.725 217.685 68.785 ;
        RECT 218.285 68.925 218.605 68.985 ;
        RECT 220.585 68.925 220.905 68.985 ;
        RECT 218.285 68.785 220.905 68.925 ;
        RECT 218.285 68.725 218.605 68.785 ;
        RECT 220.585 68.725 220.905 68.785 ;
        RECT 235.305 68.725 235.625 68.985 ;
        RECT 236.225 68.725 236.545 68.985 ;
        RECT 239.905 68.725 240.225 68.985 ;
        RECT 240.365 68.925 240.685 68.985 ;
        RECT 250.040 68.925 250.330 68.970 ;
        RECT 240.365 68.785 250.330 68.925 ;
        RECT 240.365 68.725 240.685 68.785 ;
        RECT 250.040 68.740 250.330 68.785 ;
        RECT 254.165 68.925 254.485 68.985 ;
        RECT 259.225 68.925 259.545 68.985 ;
        RECT 254.165 68.785 259.545 68.925 ;
        RECT 261.615 68.925 261.755 69.125 ;
        RECT 261.985 69.065 262.305 69.325 ;
        RECT 262.995 68.925 263.135 69.420 ;
        RECT 263.825 69.405 264.145 69.465 ;
        RECT 265.680 69.420 265.970 69.465 ;
        RECT 266.215 69.465 266.905 69.605 ;
        RECT 264.300 69.080 264.590 69.310 ;
        RECT 261.615 68.785 263.135 68.925 ;
        RECT 264.375 68.925 264.515 69.080 ;
        RECT 266.215 68.925 266.355 69.465 ;
        RECT 266.585 69.405 266.905 69.465 ;
        RECT 267.520 69.605 267.810 69.650 ;
        RECT 268.425 69.605 268.745 69.665 ;
        RECT 267.520 69.465 268.745 69.605 ;
        RECT 267.520 69.420 267.810 69.465 ;
        RECT 268.425 69.405 268.745 69.465 ;
        RECT 272.565 69.605 272.885 69.665 ;
        RECT 273.960 69.605 274.250 69.650 ;
        RECT 272.565 69.465 274.250 69.605 ;
        RECT 272.565 69.405 272.885 69.465 ;
        RECT 273.960 69.420 274.250 69.465 ;
        RECT 274.405 69.405 274.725 69.665 ;
        RECT 278.545 69.405 278.865 69.665 ;
        RECT 279.025 69.605 279.315 69.650 ;
        RECT 280.860 69.605 281.150 69.650 ;
        RECT 284.440 69.605 284.730 69.650 ;
        RECT 279.025 69.465 284.730 69.605 ;
        RECT 279.025 69.420 279.315 69.465 ;
        RECT 280.860 69.420 281.150 69.465 ;
        RECT 284.440 69.420 284.730 69.465 ;
        RECT 271.660 69.265 271.950 69.310 ;
        RECT 273.025 69.265 273.345 69.325 ;
        RECT 271.660 69.125 273.345 69.265 ;
        RECT 271.660 69.080 271.950 69.125 ;
        RECT 273.025 69.065 273.345 69.125 ;
        RECT 279.925 69.065 280.245 69.325 ;
        RECT 285.520 69.310 285.810 69.625 ;
        RECT 294.185 69.605 294.505 69.665 ;
        RECT 294.660 69.605 294.950 69.650 ;
        RECT 294.185 69.465 294.950 69.605 ;
        RECT 294.185 69.405 294.505 69.465 ;
        RECT 294.660 69.420 294.950 69.465 ;
        RECT 295.125 69.605 295.415 69.650 ;
        RECT 296.960 69.605 297.250 69.650 ;
        RECT 300.540 69.605 300.830 69.650 ;
        RECT 295.125 69.465 300.830 69.605 ;
        RECT 295.125 69.420 295.415 69.465 ;
        RECT 296.960 69.420 297.250 69.465 ;
        RECT 300.540 69.420 300.830 69.465 ;
        RECT 282.220 69.265 282.870 69.310 ;
        RECT 285.520 69.265 286.110 69.310 ;
        RECT 286.825 69.265 287.145 69.325 ;
        RECT 282.220 69.125 293.035 69.265 ;
        RECT 282.220 69.080 282.870 69.125 ;
        RECT 285.820 69.080 286.110 69.125 ;
        RECT 286.825 69.065 287.145 69.125 ;
        RECT 264.375 68.785 266.355 68.925 ;
        RECT 254.165 68.725 254.485 68.785 ;
        RECT 259.225 68.725 259.545 68.785 ;
        RECT 266.585 68.725 266.905 68.985 ;
        RECT 269.345 68.725 269.665 68.985 ;
        RECT 281.765 68.925 282.085 68.985 ;
        RECT 287.300 68.925 287.590 68.970 ;
        RECT 281.765 68.785 287.590 68.925 ;
        RECT 281.765 68.725 282.085 68.785 ;
        RECT 287.300 68.740 287.590 68.785 ;
        RECT 290.045 68.925 290.365 68.985 ;
        RECT 291.885 68.925 292.205 68.985 ;
        RECT 290.045 68.785 292.205 68.925 ;
        RECT 292.895 68.925 293.035 69.125 ;
        RECT 296.025 69.065 296.345 69.325 ;
        RECT 301.620 69.310 301.910 69.625 ;
        RECT 306.145 69.405 306.465 69.665 ;
        RECT 309.365 69.405 309.685 69.665 ;
        RECT 298.320 69.265 298.970 69.310 ;
        RECT 301.620 69.265 302.210 69.310 ;
        RECT 302.465 69.265 302.785 69.325 ;
        RECT 298.320 69.125 302.785 69.265 ;
        RECT 298.320 69.080 298.970 69.125 ;
        RECT 301.920 69.080 302.210 69.125 ;
        RECT 302.465 69.065 302.785 69.125 ;
        RECT 299.245 68.925 299.565 68.985 ;
        RECT 302.555 68.925 302.695 69.065 ;
        RECT 292.895 68.785 302.695 68.925 ;
        RECT 303.400 68.925 303.690 68.970 ;
        RECT 303.845 68.925 304.165 68.985 ;
        RECT 303.400 68.785 304.165 68.925 ;
        RECT 290.045 68.725 290.365 68.785 ;
        RECT 291.885 68.725 292.205 68.785 ;
        RECT 299.245 68.725 299.565 68.785 ;
        RECT 303.400 68.740 303.690 68.785 ;
        RECT 303.845 68.725 304.165 68.785 ;
        RECT 306.605 68.725 306.925 68.985 ;
        RECT 308.445 68.725 308.765 68.985 ;
        RECT 162.095 68.105 311.135 68.585 ;
        RECT 173.205 67.905 173.525 67.965 ;
        RECT 181.025 67.905 181.345 67.965 ;
        RECT 192.540 67.905 192.830 67.950 ;
        RECT 203.105 67.905 203.425 67.965 ;
        RECT 220.125 67.905 220.445 67.965 ;
        RECT 221.965 67.905 222.285 67.965 ;
        RECT 229.340 67.905 229.630 67.950 ;
        RECT 240.365 67.905 240.685 67.965 ;
        RECT 167.775 67.765 178.035 67.905 ;
        RECT 167.775 67.565 167.915 67.765 ;
        RECT 173.205 67.705 173.525 67.765 ;
        RECT 167.315 67.425 167.915 67.565 ;
        RECT 167.315 67.270 167.455 67.425 ;
        RECT 168.605 67.365 168.925 67.625 ;
        RECT 170.900 67.565 171.550 67.610 ;
        RECT 173.665 67.565 173.985 67.625 ;
        RECT 174.500 67.565 174.790 67.610 ;
        RECT 170.900 67.425 174.790 67.565 ;
        RECT 170.900 67.380 171.550 67.425 ;
        RECT 173.665 67.365 173.985 67.425 ;
        RECT 174.200 67.380 174.790 67.425 ;
        RECT 167.240 67.040 167.530 67.270 ;
        RECT 167.705 67.225 167.995 67.270 ;
        RECT 169.540 67.225 169.830 67.270 ;
        RECT 173.120 67.225 173.410 67.270 ;
        RECT 167.705 67.085 173.410 67.225 ;
        RECT 167.705 67.040 167.995 67.085 ;
        RECT 169.540 67.040 169.830 67.085 ;
        RECT 173.120 67.040 173.410 67.085 ;
        RECT 174.200 67.065 174.490 67.380 ;
        RECT 177.895 67.270 178.035 67.765 ;
        RECT 181.025 67.765 192.295 67.905 ;
        RECT 181.025 67.705 181.345 67.765 ;
        RECT 181.485 67.610 181.805 67.625 ;
        RECT 181.480 67.565 182.130 67.610 ;
        RECT 185.080 67.565 185.370 67.610 ;
        RECT 181.480 67.425 185.370 67.565 ;
        RECT 181.480 67.380 182.130 67.425 ;
        RECT 184.780 67.380 185.370 67.425 ;
        RECT 187.465 67.565 187.785 67.625 ;
        RECT 192.155 67.565 192.295 67.765 ;
        RECT 192.540 67.765 203.425 67.905 ;
        RECT 192.540 67.720 192.830 67.765 ;
        RECT 203.105 67.705 203.425 67.765 ;
        RECT 207.565 67.765 219.435 67.905 ;
        RECT 207.565 67.565 207.705 67.765 ;
        RECT 210.020 67.565 210.310 67.610 ;
        RECT 187.465 67.425 191.835 67.565 ;
        RECT 192.155 67.425 207.935 67.565 ;
        RECT 181.485 67.365 181.805 67.380 ;
        RECT 177.820 67.040 178.110 67.270 ;
        RECT 178.285 67.225 178.575 67.270 ;
        RECT 180.120 67.225 180.410 67.270 ;
        RECT 183.700 67.225 183.990 67.270 ;
        RECT 178.285 67.085 183.990 67.225 ;
        RECT 178.285 67.040 178.575 67.085 ;
        RECT 180.120 67.040 180.410 67.085 ;
        RECT 183.700 67.040 183.990 67.085 ;
        RECT 184.780 67.065 185.070 67.380 ;
        RECT 187.465 67.365 187.785 67.425 ;
        RECT 187.925 67.225 188.245 67.285 ;
        RECT 188.400 67.225 188.690 67.270 ;
        RECT 190.240 67.225 190.530 67.270 ;
        RECT 190.685 67.225 191.005 67.285 ;
        RECT 191.695 67.270 191.835 67.425 ;
        RECT 187.925 67.085 189.995 67.225 ;
        RECT 187.925 67.025 188.245 67.085 ;
        RECT 188.400 67.040 188.690 67.085 ;
        RECT 172.285 66.885 172.605 66.945 ;
        RECT 175.980 66.885 176.270 66.930 ;
        RECT 181.025 66.885 181.345 66.945 ;
        RECT 172.285 66.745 181.345 66.885 ;
        RECT 172.285 66.685 172.605 66.745 ;
        RECT 175.980 66.700 176.270 66.745 ;
        RECT 181.025 66.685 181.345 66.745 ;
        RECT 182.865 66.885 183.185 66.945 ;
        RECT 189.320 66.885 189.610 66.930 ;
        RECT 182.865 66.745 189.610 66.885 ;
        RECT 189.855 66.885 189.995 67.085 ;
        RECT 190.240 67.085 191.005 67.225 ;
        RECT 190.240 67.040 190.530 67.085 ;
        RECT 190.685 67.025 191.005 67.085 ;
        RECT 191.650 67.040 191.940 67.270 ;
        RECT 196.665 67.025 196.985 67.285 ;
        RECT 197.585 67.025 197.905 67.285 ;
        RECT 198.060 67.040 198.350 67.270 ;
        RECT 198.520 67.225 198.810 67.270 ;
        RECT 198.965 67.225 199.285 67.285 ;
        RECT 198.520 67.085 199.285 67.225 ;
        RECT 198.520 67.040 198.810 67.085 ;
        RECT 198.135 66.885 198.275 67.040 ;
        RECT 198.965 67.025 199.285 67.085 ;
        RECT 199.885 67.225 200.205 67.285 ;
        RECT 207.795 67.270 207.935 67.425 ;
        RECT 210.020 67.425 218.055 67.565 ;
        RECT 210.020 67.380 210.310 67.425 ;
        RECT 200.360 67.225 200.650 67.270 ;
        RECT 199.885 67.085 200.650 67.225 ;
        RECT 199.885 67.025 200.205 67.085 ;
        RECT 200.360 67.040 200.650 67.085 ;
        RECT 207.720 67.040 208.010 67.270 ;
        RECT 209.100 67.040 209.390 67.270 ;
        RECT 200.805 66.885 201.125 66.945 ;
        RECT 209.175 66.885 209.315 67.040 ;
        RECT 210.925 67.025 211.245 67.285 ;
        RECT 211.385 67.025 211.705 67.285 ;
        RECT 211.845 67.025 212.165 67.285 ;
        RECT 213.685 67.215 214.005 67.285 ;
        RECT 214.160 67.215 214.450 67.270 ;
        RECT 215.080 67.225 215.370 67.270 ;
        RECT 213.685 67.075 214.450 67.215 ;
        RECT 213.685 67.025 214.005 67.075 ;
        RECT 214.160 67.040 214.450 67.075 ;
        RECT 214.695 67.085 215.370 67.225 ;
        RECT 215.555 67.115 215.845 67.285 ;
        RECT 217.915 67.270 218.055 67.425 ;
        RECT 218.745 67.365 219.065 67.625 ;
        RECT 219.295 67.565 219.435 67.765 ;
        RECT 220.125 67.765 229.630 67.905 ;
        RECT 220.125 67.705 220.445 67.765 ;
        RECT 221.965 67.705 222.285 67.765 ;
        RECT 229.340 67.720 229.630 67.765 ;
        RECT 229.875 67.765 240.685 67.905 ;
        RECT 229.875 67.565 230.015 67.765 ;
        RECT 240.365 67.705 240.685 67.765 ;
        RECT 240.825 67.905 241.145 67.965 ;
        RECT 243.600 67.905 243.890 67.950 ;
        RECT 244.045 67.905 244.365 67.965 ;
        RECT 240.825 67.765 242.435 67.905 ;
        RECT 240.825 67.705 241.145 67.765 ;
        RECT 219.295 67.425 227.255 67.565 ;
        RECT 212.305 66.885 212.625 66.945 ;
        RECT 214.695 66.885 214.835 67.085 ;
        RECT 215.080 67.040 215.370 67.085 ;
        RECT 189.855 66.745 190.915 66.885 ;
        RECT 198.135 66.745 199.655 66.885 ;
        RECT 182.865 66.685 183.185 66.745 ;
        RECT 184.795 66.605 184.935 66.745 ;
        RECT 189.320 66.700 189.610 66.745 ;
        RECT 190.775 66.605 190.915 66.745 ;
        RECT 168.110 66.545 168.400 66.590 ;
        RECT 170.000 66.545 170.290 66.590 ;
        RECT 173.120 66.545 173.410 66.590 ;
        RECT 168.110 66.405 173.410 66.545 ;
        RECT 168.110 66.360 168.400 66.405 ;
        RECT 170.000 66.360 170.290 66.405 ;
        RECT 173.120 66.360 173.410 66.405 ;
        RECT 178.690 66.545 178.980 66.590 ;
        RECT 180.580 66.545 180.870 66.590 ;
        RECT 183.700 66.545 183.990 66.590 ;
        RECT 178.690 66.405 183.990 66.545 ;
        RECT 178.690 66.360 178.980 66.405 ;
        RECT 180.580 66.360 180.870 66.405 ;
        RECT 183.700 66.360 183.990 66.405 ;
        RECT 184.705 66.345 185.025 66.605 ;
        RECT 190.685 66.345 191.005 66.605 ;
        RECT 193.905 66.545 194.225 66.605 ;
        RECT 198.965 66.545 199.285 66.605 ;
        RECT 193.905 66.405 199.285 66.545 ;
        RECT 193.905 66.345 194.225 66.405 ;
        RECT 198.965 66.345 199.285 66.405 ;
        RECT 179.135 66.205 179.425 66.250 ;
        RECT 181.025 66.205 181.345 66.265 ;
        RECT 179.135 66.065 181.345 66.205 ;
        RECT 179.135 66.020 179.425 66.065 ;
        RECT 181.025 66.005 181.345 66.065 ;
        RECT 184.245 66.205 184.565 66.265 ;
        RECT 186.545 66.205 186.865 66.265 ;
        RECT 184.245 66.065 186.865 66.205 ;
        RECT 184.245 66.005 184.565 66.065 ;
        RECT 186.545 66.005 186.865 66.065 ;
        RECT 188.845 66.005 189.165 66.265 ;
        RECT 199.515 66.205 199.655 66.745 ;
        RECT 200.805 66.745 212.625 66.885 ;
        RECT 200.805 66.685 201.125 66.745 ;
        RECT 212.305 66.685 212.625 66.745 ;
        RECT 214.235 66.745 214.835 66.885 ;
        RECT 215.525 66.855 215.845 67.115 ;
        RECT 216.000 67.240 216.290 67.270 ;
        RECT 216.000 67.100 217.135 67.240 ;
        RECT 216.000 67.040 216.290 67.100 ;
        RECT 216.995 66.885 217.135 67.100 ;
        RECT 217.840 67.040 218.130 67.270 ;
        RECT 218.285 67.225 218.605 67.285 ;
        RECT 219.220 67.225 219.510 67.270 ;
        RECT 218.285 67.085 219.510 67.225 ;
        RECT 218.285 67.025 218.605 67.085 ;
        RECT 219.220 67.040 219.510 67.085 ;
        RECT 219.680 67.225 219.970 67.270 ;
        RECT 220.125 67.225 220.445 67.285 ;
        RECT 227.115 67.270 227.255 67.425 ;
        RECT 228.035 67.425 230.015 67.565 ;
        RECT 232.545 67.565 232.865 67.625 ;
        RECT 232.545 67.425 241.975 67.565 ;
        RECT 228.035 67.270 228.175 67.425 ;
        RECT 232.545 67.365 232.865 67.425 ;
        RECT 226.120 67.225 226.410 67.270 ;
        RECT 219.680 67.085 220.445 67.225 ;
        RECT 219.680 67.040 219.970 67.085 ;
        RECT 220.125 67.025 220.445 67.085 ;
        RECT 220.675 67.085 226.410 67.225 ;
        RECT 220.675 66.885 220.815 67.085 ;
        RECT 226.120 67.040 226.410 67.085 ;
        RECT 227.040 67.040 227.330 67.270 ;
        RECT 227.960 67.040 228.250 67.270 ;
        RECT 228.420 67.225 228.710 67.270 ;
        RECT 231.180 67.225 231.470 67.270 ;
        RECT 228.420 67.085 231.470 67.225 ;
        RECT 228.420 67.040 228.710 67.085 ;
        RECT 231.180 67.040 231.470 67.085 ;
        RECT 232.085 67.225 232.405 67.285 ;
        RECT 240.825 67.225 241.145 67.285 ;
        RECT 232.085 67.085 241.145 67.225 ;
        RECT 232.085 67.025 232.405 67.085 ;
        RECT 240.825 67.025 241.145 67.085 ;
        RECT 241.285 67.025 241.605 67.285 ;
        RECT 241.835 67.270 241.975 67.425 ;
        RECT 241.760 67.040 242.050 67.270 ;
        RECT 242.295 67.225 242.435 67.765 ;
        RECT 243.600 67.765 244.365 67.905 ;
        RECT 243.600 67.720 243.890 67.765 ;
        RECT 244.045 67.705 244.365 67.765 ;
        RECT 253.245 67.905 253.565 67.965 ;
        RECT 261.985 67.905 262.305 67.965 ;
        RECT 266.125 67.905 266.445 67.965 ;
        RECT 253.245 67.765 266.445 67.905 ;
        RECT 253.245 67.705 253.565 67.765 ;
        RECT 261.985 67.705 262.305 67.765 ;
        RECT 266.125 67.705 266.445 67.765 ;
        RECT 279.925 67.705 280.245 67.965 ;
        RECT 280.385 67.905 280.705 67.965 ;
        RECT 280.385 67.765 281.995 67.905 ;
        RECT 280.385 67.705 280.705 67.765 ;
        RECT 245.900 67.565 246.190 67.610 ;
        RECT 248.185 67.565 248.505 67.625 ;
        RECT 245.900 67.425 248.505 67.565 ;
        RECT 245.900 67.380 246.190 67.425 ;
        RECT 248.185 67.365 248.505 67.425 ;
        RECT 263.825 67.365 264.145 67.625 ;
        RECT 273.960 67.565 274.250 67.610 ;
        RECT 277.625 67.565 277.945 67.625 ;
        RECT 273.960 67.425 277.945 67.565 ;
        RECT 273.960 67.380 274.250 67.425 ;
        RECT 277.625 67.365 277.945 67.425 ;
        RECT 259.685 67.225 260.005 67.285 ;
        RECT 262.920 67.225 263.210 67.270 ;
        RECT 242.295 67.085 257.615 67.225 ;
        RECT 216.535 66.745 217.135 66.885 ;
        RECT 217.455 66.745 220.815 66.885 ;
        RECT 227.500 66.885 227.790 66.930 ;
        RECT 233.020 66.885 233.310 66.930 ;
        RECT 235.765 66.885 236.085 66.945 ;
        RECT 227.500 66.745 231.395 66.885 ;
        RECT 199.900 66.545 200.190 66.590 ;
        RECT 202.645 66.545 202.965 66.605 ;
        RECT 199.900 66.405 202.965 66.545 ;
        RECT 199.900 66.360 200.190 66.405 ;
        RECT 202.645 66.345 202.965 66.405 ;
        RECT 208.180 66.545 208.470 66.590 ;
        RECT 210.465 66.545 210.785 66.605 ;
        RECT 208.180 66.405 210.785 66.545 ;
        RECT 208.180 66.360 208.470 66.405 ;
        RECT 210.465 66.345 210.785 66.405 ;
        RECT 211.845 66.545 212.165 66.605 ;
        RECT 214.235 66.545 214.375 66.745 ;
        RECT 211.845 66.405 214.375 66.545 ;
        RECT 214.605 66.545 214.925 66.605 ;
        RECT 216.535 66.545 216.675 66.745 ;
        RECT 217.455 66.545 217.595 66.745 ;
        RECT 227.500 66.700 227.790 66.745 ;
        RECT 214.605 66.405 216.675 66.545 ;
        RECT 216.995 66.405 217.595 66.545 ;
        RECT 220.125 66.545 220.445 66.605 ;
        RECT 220.600 66.545 220.890 66.590 ;
        RECT 220.125 66.405 220.890 66.545 ;
        RECT 211.845 66.345 212.165 66.405 ;
        RECT 214.605 66.345 214.925 66.405 ;
        RECT 201.265 66.205 201.585 66.265 ;
        RECT 199.515 66.065 201.585 66.205 ;
        RECT 201.265 66.005 201.585 66.065 ;
        RECT 213.225 66.005 213.545 66.265 ;
        RECT 215.065 66.205 215.385 66.265 ;
        RECT 216.995 66.205 217.135 66.405 ;
        RECT 220.125 66.345 220.445 66.405 ;
        RECT 220.600 66.360 220.890 66.405 ;
        RECT 215.065 66.065 217.135 66.205 ;
        RECT 217.380 66.205 217.670 66.250 ;
        RECT 219.205 66.205 219.525 66.265 ;
        RECT 217.380 66.065 219.525 66.205 ;
        RECT 231.255 66.205 231.395 66.745 ;
        RECT 233.020 66.745 236.085 66.885 ;
        RECT 233.020 66.700 233.310 66.745 ;
        RECT 235.765 66.685 236.085 66.745 ;
        RECT 236.225 66.885 236.545 66.945 ;
        RECT 243.140 66.885 243.430 66.930 ;
        RECT 244.505 66.885 244.825 66.945 ;
        RECT 248.645 66.885 248.965 66.945 ;
        RECT 236.225 66.745 241.975 66.885 ;
        RECT 236.225 66.685 236.545 66.745 ;
        RECT 241.285 66.545 241.605 66.605 ;
        RECT 232.175 66.405 241.605 66.545 ;
        RECT 241.835 66.545 241.975 66.745 ;
        RECT 243.140 66.745 248.965 66.885 ;
        RECT 243.140 66.700 243.430 66.745 ;
        RECT 244.505 66.685 244.825 66.745 ;
        RECT 248.645 66.685 248.965 66.745 ;
        RECT 245.900 66.545 246.190 66.590 ;
        RECT 257.475 66.545 257.615 67.085 ;
        RECT 259.685 67.085 263.210 67.225 ;
        RECT 259.685 67.025 260.005 67.085 ;
        RECT 262.920 67.040 263.210 67.085 ;
        RECT 272.565 67.025 272.885 67.285 ;
        RECT 273.025 67.025 273.345 67.285 ;
        RECT 281.855 67.270 281.995 67.765 ;
        RECT 282.225 67.705 282.545 67.965 ;
        RECT 284.525 67.905 284.845 67.965 ;
        RECT 289.585 67.905 289.905 67.965 ;
        RECT 284.525 67.765 289.905 67.905 ;
        RECT 284.525 67.705 284.845 67.765 ;
        RECT 289.585 67.705 289.905 67.765 ;
        RECT 295.120 67.905 295.410 67.950 ;
        RECT 296.025 67.905 296.345 67.965 ;
        RECT 303.845 67.905 304.165 67.965 ;
        RECT 295.120 67.765 296.345 67.905 ;
        RECT 295.120 67.720 295.410 67.765 ;
        RECT 296.025 67.705 296.345 67.765 ;
        RECT 297.035 67.765 304.165 67.905 ;
        RECT 285.905 67.565 286.225 67.625 ;
        RECT 297.035 67.610 297.175 67.765 ;
        RECT 303.845 67.705 304.165 67.765 ;
        RECT 307.985 67.705 308.305 67.965 ;
        RECT 296.960 67.565 297.250 67.610 ;
        RECT 285.905 67.425 297.250 67.565 ;
        RECT 285.905 67.365 286.225 67.425 ;
        RECT 296.960 67.380 297.250 67.425 ;
        RECT 302.920 67.565 303.570 67.610 ;
        RECT 304.305 67.565 304.625 67.625 ;
        RECT 306.520 67.565 306.810 67.610 ;
        RECT 302.920 67.425 306.810 67.565 ;
        RECT 302.920 67.380 303.570 67.425 ;
        RECT 304.305 67.365 304.625 67.425 ;
        RECT 306.220 67.380 306.810 67.425 ;
        RECT 281.780 67.040 282.070 67.270 ;
        RECT 285.460 67.225 285.750 67.270 ;
        RECT 282.315 67.085 285.750 67.225 ;
        RECT 257.845 66.885 258.165 66.945 ;
        RECT 262.000 66.885 262.290 66.930 ;
        RECT 262.445 66.885 262.765 66.945 ;
        RECT 257.845 66.745 262.765 66.885 ;
        RECT 257.845 66.685 258.165 66.745 ;
        RECT 262.000 66.700 262.290 66.745 ;
        RECT 262.445 66.685 262.765 66.745 ;
        RECT 278.085 66.885 278.405 66.945 ;
        RECT 282.315 66.885 282.455 67.085 ;
        RECT 285.460 67.040 285.750 67.085 ;
        RECT 291.885 67.225 292.205 67.285 ;
        RECT 298.325 67.225 298.645 67.285 ;
        RECT 291.885 67.085 298.645 67.225 ;
        RECT 291.885 67.025 292.205 67.085 ;
        RECT 298.325 67.025 298.645 67.085 ;
        RECT 299.725 67.225 300.015 67.270 ;
        RECT 301.560 67.225 301.850 67.270 ;
        RECT 305.140 67.225 305.430 67.270 ;
        RECT 299.725 67.085 305.430 67.225 ;
        RECT 299.725 67.040 300.015 67.085 ;
        RECT 301.560 67.040 301.850 67.085 ;
        RECT 305.140 67.040 305.430 67.085 ;
        RECT 306.220 67.065 306.510 67.380 ;
        RECT 278.085 66.745 282.455 66.885 ;
        RECT 278.085 66.685 278.405 66.745 ;
        RECT 283.145 66.685 283.465 66.945 ;
        RECT 284.080 66.700 284.370 66.930 ;
        RECT 289.585 66.885 289.905 66.945 ;
        RECT 297.420 66.885 297.710 66.930 ;
        RECT 289.585 66.745 297.710 66.885 ;
        RECT 264.745 66.545 265.065 66.605 ;
        RECT 271.185 66.545 271.505 66.605 ;
        RECT 284.155 66.545 284.295 66.700 ;
        RECT 289.585 66.685 289.905 66.745 ;
        RECT 297.420 66.700 297.710 66.745 ;
        RECT 297.880 66.700 298.170 66.930 ;
        RECT 241.835 66.405 246.575 66.545 ;
        RECT 257.475 66.405 284.295 66.545 ;
        RECT 232.175 66.205 232.315 66.405 ;
        RECT 241.285 66.345 241.605 66.405 ;
        RECT 245.900 66.360 246.190 66.405 ;
        RECT 246.435 66.265 246.575 66.405 ;
        RECT 264.745 66.345 265.065 66.405 ;
        RECT 271.185 66.345 271.505 66.405 ;
        RECT 284.540 66.360 284.830 66.590 ;
        RECT 286.380 66.545 286.670 66.590 ;
        RECT 296.945 66.545 297.265 66.605 ;
        RECT 297.955 66.545 298.095 66.700 ;
        RECT 299.245 66.685 299.565 66.945 ;
        RECT 300.625 66.685 300.945 66.945 ;
        RECT 286.380 66.405 298.095 66.545 ;
        RECT 300.130 66.545 300.420 66.590 ;
        RECT 302.020 66.545 302.310 66.590 ;
        RECT 305.140 66.545 305.430 66.590 ;
        RECT 300.130 66.405 305.430 66.545 ;
        RECT 286.380 66.360 286.670 66.405 ;
        RECT 231.255 66.065 232.315 66.205 ;
        RECT 232.545 66.205 232.865 66.265 ;
        RECT 239.920 66.205 240.210 66.250 ;
        RECT 232.545 66.065 240.210 66.205 ;
        RECT 215.065 66.005 215.385 66.065 ;
        RECT 217.380 66.020 217.670 66.065 ;
        RECT 219.205 66.005 219.525 66.065 ;
        RECT 232.545 66.005 232.865 66.065 ;
        RECT 239.920 66.020 240.210 66.065 ;
        RECT 241.745 66.005 242.065 66.265 ;
        RECT 242.205 66.005 242.525 66.265 ;
        RECT 246.345 66.005 246.665 66.265 ;
        RECT 276.245 66.205 276.565 66.265 ;
        RECT 284.615 66.205 284.755 66.360 ;
        RECT 296.945 66.345 297.265 66.405 ;
        RECT 300.130 66.360 300.420 66.405 ;
        RECT 302.020 66.360 302.310 66.405 ;
        RECT 305.140 66.360 305.430 66.405 ;
        RECT 276.245 66.065 284.755 66.205 ;
        RECT 287.745 66.205 288.065 66.265 ;
        RECT 298.785 66.205 299.105 66.265 ;
        RECT 287.745 66.065 299.105 66.205 ;
        RECT 276.245 66.005 276.565 66.065 ;
        RECT 287.745 66.005 288.065 66.065 ;
        RECT 298.785 66.005 299.105 66.065 ;
        RECT 162.095 65.385 311.135 65.865 ;
        RECT 164.465 65.185 164.785 65.245 ;
        RECT 165.860 65.185 166.150 65.230 ;
        RECT 164.465 65.045 166.150 65.185 ;
        RECT 164.465 64.985 164.785 65.045 ;
        RECT 165.860 65.000 166.150 65.045 ;
        RECT 173.310 65.185 173.600 65.230 ;
        RECT 175.505 65.185 175.825 65.245 ;
        RECT 173.310 65.045 175.825 65.185 ;
        RECT 173.310 65.000 173.600 65.045 ;
        RECT 175.505 64.985 175.825 65.045 ;
        RECT 181.025 64.985 181.345 65.245 ;
        RECT 186.545 65.185 186.865 65.245 ;
        RECT 196.665 65.185 196.985 65.245 ;
        RECT 198.060 65.185 198.350 65.230 ;
        RECT 186.545 65.045 195.975 65.185 ;
        RECT 186.545 64.985 186.865 65.045 ;
        RECT 168.720 64.845 169.010 64.890 ;
        RECT 171.840 64.845 172.130 64.890 ;
        RECT 173.730 64.845 174.020 64.890 ;
        RECT 181.485 64.845 181.805 64.905 ;
        RECT 185.625 64.845 185.945 64.905 ;
        RECT 168.720 64.705 174.020 64.845 ;
        RECT 168.720 64.660 169.010 64.705 ;
        RECT 171.840 64.660 172.130 64.705 ;
        RECT 173.730 64.660 174.020 64.705 ;
        RECT 176.975 64.705 185.945 64.845 ;
        RECT 173.205 64.505 173.525 64.565 ;
        RECT 174.600 64.505 174.890 64.550 ;
        RECT 173.205 64.365 174.890 64.505 ;
        RECT 173.205 64.305 173.525 64.365 ;
        RECT 174.600 64.320 174.890 64.365 ;
        RECT 167.640 63.870 167.930 64.185 ;
        RECT 168.720 64.165 169.010 64.210 ;
        RECT 172.300 64.165 172.590 64.210 ;
        RECT 174.135 64.165 174.425 64.210 ;
        RECT 176.975 64.165 177.115 64.705 ;
        RECT 181.485 64.645 181.805 64.705 ;
        RECT 185.625 64.645 185.945 64.705 ;
        RECT 194.825 64.845 195.145 64.905 ;
        RECT 195.300 64.845 195.590 64.890 ;
        RECT 194.825 64.705 195.590 64.845 ;
        RECT 195.835 64.845 195.975 65.045 ;
        RECT 196.665 65.045 198.350 65.185 ;
        RECT 196.665 64.985 196.985 65.045 ;
        RECT 198.060 65.000 198.350 65.045 ;
        RECT 199.885 64.985 200.205 65.245 ;
        RECT 206.785 65.185 207.105 65.245 ;
        RECT 200.435 65.045 207.105 65.185 ;
        RECT 200.435 64.845 200.575 65.045 ;
        RECT 206.785 64.985 207.105 65.045 ;
        RECT 207.245 65.185 207.565 65.245 ;
        RECT 213.685 65.185 214.005 65.245 ;
        RECT 215.525 65.185 215.845 65.245 ;
        RECT 207.245 65.045 215.845 65.185 ;
        RECT 207.245 64.985 207.565 65.045 ;
        RECT 213.685 64.985 214.005 65.045 ;
        RECT 215.525 64.985 215.845 65.045 ;
        RECT 216.905 65.185 217.225 65.245 ;
        RECT 219.665 65.185 219.985 65.245 ;
        RECT 216.905 65.045 219.985 65.185 ;
        RECT 216.905 64.985 217.225 65.045 ;
        RECT 219.665 64.985 219.985 65.045 ;
        RECT 241.285 64.985 241.605 65.245 ;
        RECT 242.205 65.185 242.525 65.245 ;
        RECT 242.680 65.185 242.970 65.230 ;
        RECT 242.205 65.045 242.970 65.185 ;
        RECT 242.205 64.985 242.525 65.045 ;
        RECT 242.680 65.000 242.970 65.045 ;
        RECT 243.600 65.185 243.890 65.230 ;
        RECT 246.805 65.185 247.125 65.245 ;
        RECT 243.600 65.045 247.125 65.185 ;
        RECT 243.600 65.000 243.890 65.045 ;
        RECT 246.805 64.985 247.125 65.045 ;
        RECT 258.780 65.185 259.070 65.230 ;
        RECT 259.685 65.185 260.005 65.245 ;
        RECT 258.780 65.045 260.005 65.185 ;
        RECT 258.780 65.000 259.070 65.045 ;
        RECT 259.685 64.985 260.005 65.045 ;
        RECT 260.145 65.185 260.465 65.245 ;
        RECT 273.025 65.185 273.345 65.245 ;
        RECT 260.145 65.045 273.345 65.185 ;
        RECT 260.145 64.985 260.465 65.045 ;
        RECT 273.025 64.985 273.345 65.045 ;
        RECT 288.665 65.185 288.985 65.245 ;
        RECT 289.140 65.185 289.430 65.230 ;
        RECT 288.665 65.045 289.430 65.185 ;
        RECT 288.665 64.985 288.985 65.045 ;
        RECT 289.140 65.000 289.430 65.045 ;
        RECT 294.185 65.185 294.505 65.245 ;
        RECT 299.245 65.185 299.565 65.245 ;
        RECT 294.185 65.045 299.565 65.185 ;
        RECT 294.185 64.985 294.505 65.045 ;
        RECT 299.245 64.985 299.565 65.045 ;
        RECT 300.625 65.185 300.945 65.245 ;
        RECT 304.320 65.185 304.610 65.230 ;
        RECT 300.625 65.045 304.610 65.185 ;
        RECT 300.625 64.985 300.945 65.045 ;
        RECT 304.320 65.000 304.610 65.045 ;
        RECT 232.545 64.845 232.865 64.905 ;
        RECT 195.835 64.705 200.575 64.845 ;
        RECT 200.895 64.705 203.795 64.845 ;
        RECT 194.825 64.645 195.145 64.705 ;
        RECT 195.300 64.660 195.590 64.705 ;
        RECT 178.740 64.505 179.030 64.550 ;
        RECT 179.645 64.505 179.965 64.565 ;
        RECT 184.260 64.505 184.550 64.550 ;
        RECT 188.845 64.505 189.165 64.565 ;
        RECT 178.740 64.365 189.165 64.505 ;
        RECT 178.740 64.320 179.030 64.365 ;
        RECT 179.645 64.305 179.965 64.365 ;
        RECT 184.260 64.320 184.550 64.365 ;
        RECT 188.845 64.305 189.165 64.365 ;
        RECT 192.985 64.505 193.305 64.565 ;
        RECT 200.895 64.505 201.035 64.705 ;
        RECT 192.985 64.365 201.035 64.505 ;
        RECT 201.265 64.505 201.585 64.565 ;
        RECT 203.655 64.505 203.795 64.705 ;
        RECT 211.015 64.705 232.865 64.845 ;
        RECT 201.265 64.365 203.335 64.505 ;
        RECT 192.985 64.305 193.305 64.365 ;
        RECT 168.720 64.025 174.425 64.165 ;
        RECT 168.720 63.980 169.010 64.025 ;
        RECT 172.300 63.980 172.590 64.025 ;
        RECT 174.135 63.980 174.425 64.025 ;
        RECT 174.675 64.025 177.115 64.165 ;
        RECT 177.360 64.165 177.650 64.210 ;
        RECT 180.105 64.165 180.425 64.225 ;
        RECT 177.360 64.025 180.425 64.165 ;
        RECT 167.340 63.825 167.930 63.870 ;
        RECT 170.580 63.825 171.230 63.870 ;
        RECT 173.205 63.825 173.525 63.885 ;
        RECT 174.675 63.825 174.815 64.025 ;
        RECT 177.360 63.980 177.650 64.025 ;
        RECT 180.105 63.965 180.425 64.025 ;
        RECT 183.340 64.165 183.630 64.210 ;
        RECT 186.545 64.165 186.865 64.225 ;
        RECT 183.340 64.025 186.865 64.165 ;
        RECT 183.340 63.980 183.630 64.025 ;
        RECT 186.545 63.965 186.865 64.025 ;
        RECT 194.365 63.965 194.685 64.225 ;
        RECT 194.915 64.210 195.055 64.365 ;
        RECT 201.265 64.305 201.585 64.365 ;
        RECT 194.840 63.980 195.130 64.210 ;
        RECT 197.585 63.965 197.905 64.225 ;
        RECT 198.060 63.980 198.350 64.210 ;
        RECT 198.980 63.980 199.270 64.210 ;
        RECT 199.885 64.165 200.205 64.225 ;
        RECT 203.195 64.210 203.335 64.365 ;
        RECT 203.655 64.365 210.235 64.505 ;
        RECT 203.655 64.210 203.795 64.365 ;
        RECT 202.660 64.165 202.950 64.210 ;
        RECT 199.885 64.025 202.950 64.165 ;
        RECT 177.820 63.825 178.110 63.870 ;
        RECT 193.905 63.825 194.225 63.885 ;
        RECT 167.340 63.685 174.815 63.825 ;
        RECT 175.135 63.685 194.225 63.825 ;
        RECT 167.340 63.640 167.630 63.685 ;
        RECT 170.580 63.640 171.230 63.685 ;
        RECT 173.205 63.625 173.525 63.685 ;
        RECT 169.065 63.485 169.385 63.545 ;
        RECT 175.135 63.485 175.275 63.685 ;
        RECT 177.820 63.640 178.110 63.685 ;
        RECT 193.905 63.625 194.225 63.685 ;
        RECT 195.745 63.825 196.065 63.885 ;
        RECT 198.135 63.825 198.275 63.980 ;
        RECT 195.745 63.685 198.275 63.825 ;
        RECT 199.055 63.825 199.195 63.980 ;
        RECT 199.885 63.965 200.205 64.025 ;
        RECT 202.660 63.980 202.950 64.025 ;
        RECT 203.120 63.980 203.410 64.210 ;
        RECT 203.580 63.980 203.870 64.210 ;
        RECT 200.345 63.825 200.665 63.885 ;
        RECT 199.055 63.685 200.665 63.825 ;
        RECT 203.195 63.825 203.335 63.980 ;
        RECT 204.485 63.965 204.805 64.225 ;
        RECT 207.245 63.965 207.565 64.225 ;
        RECT 208.180 63.980 208.470 64.210 ;
        RECT 208.255 63.825 208.395 63.980 ;
        RECT 208.625 63.965 208.945 64.225 ;
        RECT 209.100 64.165 209.390 64.210 ;
        RECT 209.545 64.165 209.865 64.225 ;
        RECT 209.100 64.025 209.865 64.165 ;
        RECT 210.095 64.165 210.235 64.365 ;
        RECT 210.465 64.305 210.785 64.565 ;
        RECT 211.015 64.210 211.155 64.705 ;
        RECT 210.095 64.025 210.695 64.165 ;
        RECT 209.100 63.980 209.390 64.025 ;
        RECT 209.545 63.965 209.865 64.025 ;
        RECT 210.005 63.825 210.325 63.885 ;
        RECT 203.195 63.685 207.705 63.825 ;
        RECT 208.255 63.685 210.325 63.825 ;
        RECT 210.555 63.825 210.695 64.025 ;
        RECT 210.940 63.980 211.230 64.210 ;
        RECT 211.845 63.965 212.165 64.225 ;
        RECT 212.320 63.980 212.610 64.210 ;
        RECT 211.935 63.825 212.075 63.965 ;
        RECT 210.555 63.685 212.075 63.825 ;
        RECT 195.745 63.625 196.065 63.685 ;
        RECT 200.345 63.625 200.665 63.685 ;
        RECT 169.065 63.345 175.275 63.485 ;
        RECT 175.520 63.485 175.810 63.530 ;
        RECT 175.965 63.485 176.285 63.545 ;
        RECT 175.520 63.345 176.285 63.485 ;
        RECT 169.065 63.285 169.385 63.345 ;
        RECT 175.520 63.300 175.810 63.345 ;
        RECT 175.965 63.285 176.285 63.345 ;
        RECT 182.880 63.485 183.170 63.530 ;
        RECT 190.225 63.485 190.545 63.545 ;
        RECT 182.880 63.345 190.545 63.485 ;
        RECT 182.880 63.300 183.170 63.345 ;
        RECT 190.225 63.285 190.545 63.345 ;
        RECT 198.965 63.485 199.285 63.545 ;
        RECT 201.280 63.485 201.570 63.530 ;
        RECT 198.965 63.345 201.570 63.485 ;
        RECT 207.565 63.485 207.705 63.685 ;
        RECT 210.005 63.625 210.325 63.685 ;
        RECT 208.625 63.485 208.945 63.545 ;
        RECT 212.395 63.485 212.535 63.980 ;
        RECT 212.765 63.965 213.085 64.225 ;
        RECT 214.650 64.175 214.940 64.210 ;
        RECT 215.155 64.175 215.295 64.705 ;
        RECT 232.545 64.645 232.865 64.705 ;
        RECT 244.045 64.845 244.365 64.905 ;
        RECT 263.365 64.845 263.685 64.905 ;
        RECT 279.465 64.845 279.785 64.905 ;
        RECT 244.045 64.705 279.785 64.845 ;
        RECT 244.045 64.645 244.365 64.705 ;
        RECT 263.365 64.645 263.685 64.705 ;
        RECT 279.465 64.645 279.785 64.705 ;
        RECT 281.270 64.845 281.560 64.890 ;
        RECT 283.160 64.845 283.450 64.890 ;
        RECT 286.280 64.845 286.570 64.890 ;
        RECT 281.270 64.705 286.570 64.845 ;
        RECT 281.270 64.660 281.560 64.705 ;
        RECT 283.160 64.660 283.450 64.705 ;
        RECT 286.280 64.660 286.570 64.705 ;
        RECT 295.070 64.845 295.360 64.890 ;
        RECT 296.960 64.845 297.250 64.890 ;
        RECT 300.080 64.845 300.370 64.890 ;
        RECT 295.070 64.705 300.370 64.845 ;
        RECT 295.070 64.660 295.360 64.705 ;
        RECT 296.960 64.660 297.250 64.705 ;
        RECT 300.080 64.660 300.370 64.705 ;
        RECT 218.745 64.505 219.065 64.565 ;
        RECT 220.140 64.505 220.430 64.550 ;
        RECT 218.745 64.365 220.430 64.505 ;
        RECT 218.745 64.305 219.065 64.365 ;
        RECT 220.140 64.320 220.430 64.365 ;
        RECT 221.045 64.505 221.365 64.565 ;
        RECT 278.085 64.505 278.405 64.565 ;
        RECT 221.045 64.365 278.405 64.505 ;
        RECT 221.045 64.305 221.365 64.365 ;
        RECT 214.650 64.035 215.295 64.175 ;
        RECT 214.650 63.980 214.940 64.035 ;
        RECT 215.525 63.965 215.845 64.225 ;
        RECT 216.000 63.980 216.290 64.210 ;
        RECT 216.460 64.165 216.750 64.210 ;
        RECT 216.905 64.165 217.225 64.225 ;
        RECT 216.460 64.025 217.225 64.165 ;
        RECT 216.460 63.980 216.750 64.025 ;
        RECT 213.685 63.825 214.005 63.885 ;
        RECT 214.160 63.825 214.450 63.870 ;
        RECT 213.685 63.685 214.450 63.825 ;
        RECT 213.685 63.625 214.005 63.685 ;
        RECT 214.160 63.640 214.450 63.685 ;
        RECT 215.065 63.825 215.385 63.885 ;
        RECT 216.075 63.825 216.215 63.980 ;
        RECT 216.905 63.965 217.225 64.025 ;
        RECT 219.205 63.965 219.525 64.225 ;
        RECT 219.665 63.965 219.985 64.225 ;
        RECT 220.585 63.965 220.905 64.225 ;
        RECT 221.520 64.165 221.810 64.210 ;
        RECT 225.185 64.165 225.505 64.225 ;
        RECT 221.520 64.025 225.505 64.165 ;
        RECT 221.520 63.980 221.810 64.025 ;
        RECT 225.185 63.965 225.505 64.025 ;
        RECT 243.125 63.965 243.445 64.225 ;
        RECT 244.060 64.165 244.350 64.210 ;
        RECT 244.505 64.165 244.825 64.225 ;
        RECT 244.060 64.025 244.825 64.165 ;
        RECT 244.060 63.980 244.350 64.025 ;
        RECT 244.505 63.965 244.825 64.025 ;
        RECT 244.980 64.165 245.270 64.210 ;
        RECT 247.265 64.165 247.585 64.225 ;
        RECT 244.980 64.025 247.585 64.165 ;
        RECT 244.980 63.980 245.270 64.025 ;
        RECT 247.265 63.965 247.585 64.025 ;
        RECT 256.925 63.965 257.245 64.225 ;
        RECT 257.935 64.210 258.075 64.365 ;
        RECT 278.085 64.305 278.405 64.365 ;
        RECT 278.545 64.505 278.865 64.565 ;
        RECT 280.400 64.505 280.690 64.550 ;
        RECT 294.185 64.505 294.505 64.565 ;
        RECT 278.545 64.365 294.505 64.505 ;
        RECT 278.545 64.305 278.865 64.365 ;
        RECT 280.400 64.320 280.690 64.365 ;
        RECT 294.185 64.305 294.505 64.365 ;
        RECT 297.405 64.505 297.725 64.565 ;
        RECT 307.080 64.505 307.370 64.550 ;
        RECT 297.405 64.365 307.370 64.505 ;
        RECT 297.405 64.305 297.725 64.365 ;
        RECT 307.080 64.320 307.370 64.365 ;
        RECT 257.860 63.980 258.150 64.210 ;
        RECT 259.240 64.165 259.530 64.210 ;
        RECT 276.245 64.165 276.565 64.225 ;
        RECT 259.240 64.025 276.565 64.165 ;
        RECT 259.240 63.980 259.530 64.025 ;
        RECT 215.065 63.685 216.215 63.825 ;
        RECT 217.840 63.825 218.130 63.870 ;
        RECT 226.105 63.825 226.425 63.885 ;
        RECT 217.840 63.685 226.425 63.825 ;
        RECT 215.065 63.625 215.385 63.685 ;
        RECT 217.840 63.640 218.130 63.685 ;
        RECT 226.105 63.625 226.425 63.685 ;
        RECT 231.625 63.825 231.945 63.885 ;
        RECT 259.315 63.825 259.455 63.980 ;
        RECT 276.245 63.965 276.565 64.025 ;
        RECT 280.865 64.165 281.155 64.210 ;
        RECT 282.700 64.165 282.990 64.210 ;
        RECT 286.280 64.165 286.570 64.210 ;
        RECT 280.865 64.025 286.570 64.165 ;
        RECT 280.865 63.980 281.155 64.025 ;
        RECT 282.700 63.980 282.990 64.025 ;
        RECT 286.280 63.980 286.570 64.025 ;
        RECT 231.625 63.685 259.455 63.825 ;
        RECT 260.605 63.825 260.925 63.885 ;
        RECT 272.120 63.825 272.410 63.870 ;
        RECT 272.565 63.825 272.885 63.885 ;
        RECT 260.605 63.685 272.885 63.825 ;
        RECT 231.625 63.625 231.945 63.685 ;
        RECT 260.605 63.625 260.925 63.685 ;
        RECT 272.120 63.640 272.410 63.685 ;
        RECT 272.565 63.625 272.885 63.685 ;
        RECT 273.040 63.825 273.330 63.870 ;
        RECT 274.405 63.825 274.725 63.885 ;
        RECT 273.040 63.685 274.725 63.825 ;
        RECT 273.040 63.640 273.330 63.685 ;
        RECT 274.405 63.625 274.725 63.685 ;
        RECT 281.780 63.825 282.070 63.870 ;
        RECT 282.225 63.825 282.545 63.885 ;
        RECT 281.780 63.685 282.545 63.825 ;
        RECT 281.780 63.640 282.070 63.685 ;
        RECT 282.225 63.625 282.545 63.685 ;
        RECT 284.060 63.825 284.710 63.870 ;
        RECT 286.825 63.825 287.145 63.885 ;
        RECT 287.360 63.870 287.650 64.185 ;
        RECT 294.665 64.165 294.955 64.210 ;
        RECT 296.500 64.165 296.790 64.210 ;
        RECT 300.080 64.165 300.370 64.210 ;
        RECT 294.665 64.025 300.370 64.165 ;
        RECT 294.665 63.980 294.955 64.025 ;
        RECT 296.500 63.980 296.790 64.025 ;
        RECT 300.080 63.980 300.370 64.025 ;
        RECT 287.360 63.825 287.950 63.870 ;
        RECT 284.060 63.685 287.950 63.825 ;
        RECT 284.060 63.640 284.710 63.685 ;
        RECT 286.825 63.625 287.145 63.685 ;
        RECT 287.660 63.640 287.950 63.685 ;
        RECT 295.105 63.825 295.425 63.885 ;
        RECT 297.865 63.870 298.185 63.885 ;
        RECT 301.160 63.870 301.450 64.185 ;
        RECT 306.160 64.165 306.450 64.210 ;
        RECT 307.985 64.165 308.305 64.225 ;
        RECT 306.160 64.025 308.305 64.165 ;
        RECT 306.160 63.980 306.450 64.025 ;
        RECT 307.985 63.965 308.305 64.025 ;
        RECT 295.580 63.825 295.870 63.870 ;
        RECT 295.105 63.685 295.870 63.825 ;
        RECT 295.105 63.625 295.425 63.685 ;
        RECT 295.580 63.640 295.870 63.685 ;
        RECT 297.860 63.825 298.510 63.870 ;
        RECT 301.160 63.825 301.750 63.870 ;
        RECT 297.860 63.685 301.750 63.825 ;
        RECT 297.860 63.640 298.510 63.685 ;
        RECT 301.460 63.640 301.750 63.685 ;
        RECT 297.865 63.625 298.185 63.640 ;
        RECT 215.155 63.485 215.295 63.625 ;
        RECT 207.565 63.345 215.295 63.485 ;
        RECT 198.965 63.285 199.285 63.345 ;
        RECT 201.280 63.300 201.570 63.345 ;
        RECT 208.625 63.285 208.945 63.345 ;
        RECT 218.285 63.285 218.605 63.545 ;
        RECT 231.165 63.485 231.485 63.545 ;
        RECT 270.725 63.485 271.045 63.545 ;
        RECT 231.165 63.345 271.045 63.485 ;
        RECT 231.165 63.285 231.485 63.345 ;
        RECT 270.725 63.285 271.045 63.345 ;
        RECT 271.185 63.485 271.505 63.545 ;
        RECT 273.960 63.485 274.250 63.530 ;
        RECT 271.185 63.345 274.250 63.485 ;
        RECT 271.185 63.285 271.505 63.345 ;
        RECT 273.960 63.300 274.250 63.345 ;
        RECT 281.305 63.485 281.625 63.545 ;
        RECT 290.045 63.485 290.365 63.545 ;
        RECT 281.305 63.345 290.365 63.485 ;
        RECT 281.305 63.285 281.625 63.345 ;
        RECT 290.045 63.285 290.365 63.345 ;
        RECT 296.485 63.485 296.805 63.545 ;
        RECT 302.940 63.485 303.230 63.530 ;
        RECT 305.685 63.485 306.005 63.545 ;
        RECT 296.485 63.345 306.005 63.485 ;
        RECT 296.485 63.285 296.805 63.345 ;
        RECT 302.940 63.300 303.230 63.345 ;
        RECT 305.685 63.285 306.005 63.345 ;
        RECT 306.605 63.285 306.925 63.545 ;
        RECT 162.095 62.665 311.135 63.145 ;
        RECT 168.620 62.465 168.910 62.510 ;
        RECT 169.065 62.465 169.385 62.525 ;
        RECT 168.620 62.325 169.385 62.465 ;
        RECT 168.620 62.280 168.910 62.325 ;
        RECT 169.065 62.265 169.385 62.325 ;
        RECT 178.280 62.465 178.570 62.510 ;
        RECT 180.105 62.465 180.425 62.525 ;
        RECT 178.280 62.325 180.425 62.465 ;
        RECT 178.280 62.280 178.570 62.325 ;
        RECT 180.105 62.265 180.425 62.325 ;
        RECT 186.100 62.465 186.390 62.510 ;
        RECT 188.385 62.465 188.705 62.525 ;
        RECT 186.100 62.325 188.705 62.465 ;
        RECT 186.100 62.280 186.390 62.325 ;
        RECT 188.385 62.265 188.705 62.325 ;
        RECT 189.305 62.265 189.625 62.525 ;
        RECT 190.700 62.465 190.990 62.510 ;
        RECT 191.145 62.465 191.465 62.525 ;
        RECT 190.700 62.325 191.465 62.465 ;
        RECT 190.700 62.280 190.990 62.325 ;
        RECT 191.145 62.265 191.465 62.325 ;
        RECT 194.840 62.465 195.130 62.510 ;
        RECT 197.125 62.465 197.445 62.525 ;
        RECT 194.840 62.325 197.445 62.465 ;
        RECT 194.840 62.280 195.130 62.325 ;
        RECT 197.125 62.265 197.445 62.325 ;
        RECT 197.585 62.465 197.905 62.525 ;
        RECT 202.200 62.465 202.490 62.510 ;
        RECT 207.245 62.465 207.565 62.525 ;
        RECT 197.585 62.325 207.565 62.465 ;
        RECT 197.585 62.265 197.905 62.325 ;
        RECT 202.200 62.280 202.490 62.325 ;
        RECT 207.245 62.265 207.565 62.325 ;
        RECT 208.165 62.465 208.485 62.525 ;
        RECT 221.045 62.465 221.365 62.525 ;
        RECT 208.165 62.325 221.365 62.465 ;
        RECT 208.165 62.265 208.485 62.325 ;
        RECT 221.045 62.265 221.365 62.325 ;
        RECT 231.165 62.265 231.485 62.525 ;
        RECT 234.860 62.465 235.150 62.510 ;
        RECT 239.445 62.465 239.765 62.525 ;
        RECT 241.300 62.465 241.590 62.510 ;
        RECT 234.860 62.325 241.590 62.465 ;
        RECT 234.860 62.280 235.150 62.325 ;
        RECT 239.445 62.265 239.765 62.325 ;
        RECT 241.300 62.280 241.590 62.325 ;
        RECT 241.760 62.465 242.050 62.510 ;
        RECT 242.205 62.465 242.525 62.525 ;
        RECT 241.760 62.325 242.525 62.465 ;
        RECT 241.760 62.280 242.050 62.325 ;
        RECT 242.205 62.265 242.525 62.325 ;
        RECT 243.125 62.265 243.445 62.525 ;
        RECT 243.585 62.465 243.905 62.525 ;
        RECT 244.520 62.465 244.810 62.510 ;
        RECT 248.185 62.465 248.505 62.525 ;
        RECT 243.585 62.325 248.505 62.465 ;
        RECT 243.585 62.265 243.905 62.325 ;
        RECT 244.520 62.280 244.810 62.325 ;
        RECT 248.185 62.265 248.505 62.325 ;
        RECT 252.325 62.465 252.645 62.525 ;
        RECT 255.545 62.465 255.865 62.525 ;
        RECT 252.325 62.325 255.865 62.465 ;
        RECT 252.325 62.265 252.645 62.325 ;
        RECT 255.545 62.265 255.865 62.325 ;
        RECT 256.940 62.465 257.230 62.510 ;
        RECT 257.845 62.465 258.165 62.525 ;
        RECT 260.605 62.510 260.925 62.525 ;
        RECT 260.575 62.465 260.925 62.510 ;
        RECT 256.940 62.325 258.165 62.465 ;
        RECT 260.410 62.325 260.925 62.465 ;
        RECT 256.940 62.280 257.230 62.325 ;
        RECT 257.845 62.265 258.165 62.325 ;
        RECT 260.575 62.280 260.925 62.325 ;
        RECT 260.605 62.265 260.925 62.280 ;
        RECT 270.725 62.465 271.045 62.525 ;
        RECT 280.845 62.465 281.165 62.525 ;
        RECT 270.725 62.325 281.995 62.465 ;
        RECT 270.725 62.265 271.045 62.325 ;
        RECT 280.845 62.265 281.165 62.325 ;
        RECT 173.205 62.170 173.525 62.185 ;
        RECT 170.100 62.125 170.390 62.170 ;
        RECT 173.205 62.125 173.990 62.170 ;
        RECT 170.100 61.985 173.990 62.125 ;
        RECT 170.100 61.940 170.690 61.985 ;
        RECT 164.925 61.585 165.245 61.845 ;
        RECT 170.400 61.625 170.690 61.940 ;
        RECT 173.205 61.940 173.990 61.985 ;
        RECT 173.205 61.925 173.525 61.940 ;
        RECT 175.965 61.925 176.285 62.185 ;
        RECT 189.395 62.125 189.535 62.265 ;
        RECT 180.195 61.985 189.535 62.125 ;
        RECT 194.365 62.125 194.685 62.185 ;
        RECT 220.585 62.125 220.905 62.185 ;
        RECT 224.740 62.125 225.030 62.170 ;
        RECT 247.725 62.125 248.045 62.185 ;
        RECT 194.365 61.985 201.495 62.125 ;
        RECT 180.195 61.845 180.335 61.985 ;
        RECT 194.365 61.925 194.685 61.985 ;
        RECT 171.480 61.785 171.770 61.830 ;
        RECT 175.060 61.785 175.350 61.830 ;
        RECT 176.895 61.785 177.185 61.830 ;
        RECT 171.480 61.645 177.185 61.785 ;
        RECT 171.480 61.600 171.770 61.645 ;
        RECT 175.060 61.600 175.350 61.645 ;
        RECT 176.895 61.600 177.185 61.645 ;
        RECT 179.200 61.785 179.490 61.830 ;
        RECT 179.645 61.785 179.965 61.845 ;
        RECT 179.200 61.645 179.965 61.785 ;
        RECT 179.200 61.600 179.490 61.645 ;
        RECT 179.645 61.585 179.965 61.645 ;
        RECT 180.105 61.585 180.425 61.845 ;
        RECT 184.245 61.785 184.565 61.845 ;
        RECT 186.100 61.785 186.390 61.830 ;
        RECT 184.245 61.645 186.390 61.785 ;
        RECT 184.245 61.585 184.565 61.645 ;
        RECT 186.100 61.600 186.390 61.645 ;
        RECT 188.385 61.585 188.705 61.845 ;
        RECT 189.305 61.785 189.625 61.845 ;
        RECT 192.540 61.785 192.830 61.830 ;
        RECT 189.305 61.645 192.830 61.785 ;
        RECT 189.305 61.585 189.625 61.645 ;
        RECT 192.540 61.600 192.830 61.645 ;
        RECT 177.360 61.260 177.650 61.490 ;
        RECT 171.480 61.105 171.770 61.150 ;
        RECT 174.600 61.105 174.890 61.150 ;
        RECT 176.490 61.105 176.780 61.150 ;
        RECT 171.480 60.965 176.780 61.105 ;
        RECT 171.480 60.920 171.770 60.965 ;
        RECT 174.600 60.920 174.890 60.965 ;
        RECT 176.490 60.920 176.780 60.965 ;
        RECT 164.005 60.565 164.325 60.825 ;
        RECT 175.045 60.765 175.365 60.825 ;
        RECT 177.435 60.765 177.575 61.260 ;
        RECT 184.705 61.245 185.025 61.505 ;
        RECT 187.465 61.445 187.785 61.505 ;
        RECT 189.780 61.445 190.070 61.490 ;
        RECT 187.465 61.305 190.070 61.445 ;
        RECT 187.465 61.245 187.785 61.305 ;
        RECT 189.780 61.260 190.070 61.305 ;
        RECT 185.640 60.920 185.930 61.150 ;
        RECT 175.045 60.625 177.575 60.765 ;
        RECT 185.715 60.765 185.855 60.920 ;
        RECT 188.845 60.905 189.165 61.165 ;
        RECT 194.380 61.105 194.670 61.150 ;
        RECT 194.915 61.105 195.055 61.985 ;
        RECT 197.600 61.600 197.890 61.830 ;
        RECT 197.675 61.445 197.815 61.600 ;
        RECT 198.045 61.585 198.365 61.845 ;
        RECT 198.505 61.585 198.825 61.845 ;
        RECT 198.965 61.585 199.285 61.845 ;
        RECT 199.885 61.585 200.205 61.845 ;
        RECT 200.345 61.585 200.665 61.845 ;
        RECT 201.355 61.830 201.495 61.985 ;
        RECT 211.015 61.985 218.055 62.125 ;
        RECT 211.015 61.845 211.155 61.985 ;
        RECT 201.280 61.600 201.570 61.830 ;
        RECT 208.625 61.585 208.945 61.845 ;
        RECT 209.085 61.785 209.405 61.845 ;
        RECT 209.560 61.785 209.850 61.830 ;
        RECT 209.085 61.645 209.850 61.785 ;
        RECT 209.085 61.585 209.405 61.645 ;
        RECT 209.560 61.600 209.850 61.645 ;
        RECT 210.925 61.585 211.245 61.845 ;
        RECT 212.305 61.585 212.625 61.845 ;
        RECT 215.525 61.585 215.845 61.845 ;
        RECT 215.985 61.585 216.305 61.845 ;
        RECT 216.445 61.585 216.765 61.845 ;
        RECT 217.915 61.830 218.055 61.985 ;
        RECT 220.585 61.985 248.045 62.125 ;
        RECT 248.275 62.125 248.415 62.265 ;
        RECT 262.460 62.125 262.750 62.170 ;
        RECT 274.405 62.125 274.725 62.185 ;
        RECT 248.275 61.985 274.725 62.125 ;
        RECT 220.585 61.925 220.905 61.985 ;
        RECT 224.740 61.940 225.030 61.985 ;
        RECT 247.725 61.925 248.045 61.985 ;
        RECT 262.460 61.940 262.750 61.985 ;
        RECT 274.405 61.925 274.725 61.985 ;
        RECT 278.085 62.125 278.405 62.185 ;
        RECT 278.085 61.985 281.075 62.125 ;
        RECT 278.085 61.925 278.405 61.985 ;
        RECT 217.840 61.785 218.130 61.830 ;
        RECT 226.120 61.785 226.410 61.830 ;
        RECT 217.840 61.645 226.410 61.785 ;
        RECT 217.840 61.600 218.130 61.645 ;
        RECT 226.120 61.600 226.410 61.645 ;
        RECT 226.565 61.785 226.885 61.845 ;
        RECT 227.040 61.785 227.330 61.830 ;
        RECT 226.565 61.645 227.330 61.785 ;
        RECT 226.565 61.585 226.885 61.645 ;
        RECT 227.040 61.600 227.330 61.645 ;
        RECT 227.500 61.600 227.790 61.830 ;
        RECT 203.105 61.445 203.425 61.505 ;
        RECT 197.675 61.305 203.425 61.445 ;
        RECT 203.105 61.245 203.425 61.305 ;
        RECT 211.845 61.445 212.165 61.505 ;
        RECT 213.240 61.445 213.530 61.490 ;
        RECT 211.845 61.305 213.530 61.445 ;
        RECT 211.845 61.245 212.165 61.305 ;
        RECT 213.240 61.260 213.530 61.305 ;
        RECT 213.685 61.445 214.005 61.505 ;
        RECT 216.920 61.445 217.210 61.490 ;
        RECT 213.685 61.305 217.210 61.445 ;
        RECT 213.685 61.245 214.005 61.305 ;
        RECT 216.920 61.260 217.210 61.305 ;
        RECT 221.505 61.245 221.825 61.505 ;
        RECT 227.575 61.445 227.715 61.600 ;
        RECT 230.705 61.585 231.025 61.845 ;
        RECT 234.845 61.785 235.165 61.845 ;
        RECT 235.320 61.785 235.610 61.830 ;
        RECT 234.845 61.645 235.610 61.785 ;
        RECT 234.845 61.585 235.165 61.645 ;
        RECT 235.320 61.600 235.610 61.645 ;
        RECT 236.685 61.785 237.005 61.845 ;
        RECT 239.920 61.785 240.210 61.830 ;
        RECT 243.585 61.785 243.905 61.845 ;
        RECT 236.685 61.645 243.905 61.785 ;
        RECT 236.685 61.585 237.005 61.645 ;
        RECT 239.920 61.600 240.210 61.645 ;
        RECT 243.585 61.585 243.905 61.645 ;
        RECT 244.045 61.585 244.365 61.845 ;
        RECT 244.505 61.785 244.825 61.845 ;
        RECT 245.440 61.785 245.730 61.830 ;
        RECT 244.505 61.645 245.730 61.785 ;
        RECT 244.505 61.585 244.825 61.645 ;
        RECT 245.440 61.600 245.730 61.645 ;
        RECT 246.805 61.585 247.125 61.845 ;
        RECT 252.785 61.585 253.105 61.845 ;
        RECT 259.240 61.785 259.530 61.830 ;
        RECT 259.685 61.785 260.005 61.845 ;
        RECT 259.240 61.645 260.005 61.785 ;
        RECT 259.240 61.600 259.530 61.645 ;
        RECT 259.685 61.585 260.005 61.645 ;
        RECT 276.245 61.785 276.565 61.845 ;
        RECT 280.935 61.830 281.075 61.985 ;
        RECT 279.480 61.785 279.770 61.830 ;
        RECT 276.245 61.645 279.770 61.785 ;
        RECT 276.245 61.585 276.565 61.645 ;
        RECT 279.480 61.600 279.770 61.645 ;
        RECT 280.860 61.600 281.150 61.830 ;
        RECT 281.855 61.785 281.995 62.325 ;
        RECT 282.225 62.265 282.545 62.525 ;
        RECT 284.080 62.465 284.370 62.510 ;
        RECT 288.665 62.465 288.985 62.525 ;
        RECT 284.080 62.325 288.985 62.465 ;
        RECT 284.080 62.280 284.370 62.325 ;
        RECT 288.665 62.265 288.985 62.325 ;
        RECT 295.105 62.265 295.425 62.525 ;
        RECT 296.025 62.465 296.345 62.525 ;
        RECT 297.420 62.465 297.710 62.510 ;
        RECT 306.605 62.465 306.925 62.525 ;
        RECT 296.025 62.325 297.710 62.465 ;
        RECT 296.025 62.265 296.345 62.325 ;
        RECT 297.420 62.280 297.710 62.325 ;
        RECT 300.715 62.325 306.925 62.465 ;
        RECT 296.485 62.125 296.805 62.185 ;
        RECT 296.960 62.125 297.250 62.170 ;
        RECT 296.485 61.985 297.250 62.125 ;
        RECT 296.485 61.925 296.805 61.985 ;
        RECT 296.960 61.940 297.250 61.985 ;
        RECT 287.745 61.785 288.065 61.845 ;
        RECT 288.220 61.785 288.510 61.830 ;
        RECT 300.715 61.785 300.855 62.325 ;
        RECT 306.605 62.265 306.925 62.325 ;
        RECT 302.465 62.125 302.785 62.185 ;
        RECT 303.400 62.125 303.690 62.170 ;
        RECT 302.465 61.985 303.690 62.125 ;
        RECT 302.465 61.925 302.785 61.985 ;
        RECT 303.400 61.940 303.690 61.985 ;
        RECT 305.225 61.925 305.545 62.185 ;
        RECT 281.855 61.645 287.515 61.785 ;
        RECT 224.355 61.305 227.715 61.445 ;
        RECT 232.100 61.445 232.390 61.490 ;
        RECT 235.780 61.445 236.070 61.490 ;
        RECT 232.100 61.305 236.070 61.445 ;
        RECT 200.345 61.105 200.665 61.165 ;
        RECT 194.380 60.965 195.055 61.105 ;
        RECT 195.375 60.965 200.665 61.105 ;
        RECT 194.380 60.920 194.670 60.965 ;
        RECT 186.085 60.765 186.405 60.825 ;
        RECT 191.605 60.765 191.925 60.825 ;
        RECT 195.375 60.765 195.515 60.965 ;
        RECT 200.345 60.905 200.665 60.965 ;
        RECT 207.705 61.105 208.025 61.165 ;
        RECT 209.100 61.105 209.390 61.150 ;
        RECT 207.705 60.965 209.390 61.105 ;
        RECT 207.705 60.905 208.025 60.965 ;
        RECT 209.100 60.920 209.390 60.965 ;
        RECT 221.045 61.105 221.365 61.165 ;
        RECT 224.355 61.105 224.495 61.305 ;
        RECT 232.100 61.260 232.390 61.305 ;
        RECT 235.780 61.260 236.070 61.305 ;
        RECT 242.345 61.445 242.635 61.490 ;
        RECT 246.345 61.445 246.665 61.505 ;
        RECT 242.345 61.305 246.665 61.445 ;
        RECT 242.345 61.260 242.635 61.305 ;
        RECT 221.045 60.965 224.495 61.105 ;
        RECT 226.105 61.105 226.425 61.165 ;
        RECT 226.580 61.105 226.870 61.150 ;
        RECT 226.105 60.965 226.870 61.105 ;
        RECT 235.855 61.105 235.995 61.260 ;
        RECT 246.345 61.245 246.665 61.305 ;
        RECT 251.420 61.260 251.710 61.490 ;
        RECT 251.495 61.105 251.635 61.260 ;
        RECT 257.385 61.245 257.705 61.505 ;
        RECT 257.860 61.260 258.150 61.490 ;
        RECT 279.925 61.445 280.245 61.505 ;
        RECT 282.685 61.445 283.005 61.505 ;
        RECT 258.395 61.305 269.805 61.445 ;
        RECT 256.925 61.105 257.245 61.165 ;
        RECT 257.935 61.105 258.075 61.260 ;
        RECT 235.855 60.965 258.075 61.105 ;
        RECT 221.045 60.905 221.365 60.965 ;
        RECT 226.105 60.905 226.425 60.965 ;
        RECT 226.580 60.920 226.870 60.965 ;
        RECT 256.925 60.905 257.245 60.965 ;
        RECT 185.715 60.625 195.515 60.765 ;
        RECT 175.045 60.565 175.365 60.625 ;
        RECT 186.085 60.565 186.405 60.625 ;
        RECT 191.605 60.565 191.925 60.625 ;
        RECT 196.205 60.565 196.525 60.825 ;
        RECT 207.245 60.565 207.565 60.825 ;
        RECT 210.020 60.765 210.310 60.810 ;
        RECT 211.400 60.765 211.690 60.810 ;
        RECT 210.020 60.625 211.690 60.765 ;
        RECT 210.020 60.580 210.310 60.625 ;
        RECT 211.400 60.580 211.690 60.625 ;
        RECT 211.845 60.765 212.165 60.825 ;
        RECT 214.160 60.765 214.450 60.810 ;
        RECT 211.845 60.625 214.450 60.765 ;
        RECT 211.845 60.565 212.165 60.625 ;
        RECT 214.160 60.580 214.450 60.625 ;
        RECT 225.185 60.565 225.505 60.825 ;
        RECT 228.865 60.565 229.185 60.825 ;
        RECT 232.545 60.765 232.865 60.825 ;
        RECT 233.020 60.765 233.310 60.810 ;
        RECT 232.545 60.625 233.310 60.765 ;
        RECT 232.545 60.565 232.865 60.625 ;
        RECT 233.020 60.580 233.310 60.625 ;
        RECT 246.345 60.565 246.665 60.825 ;
        RECT 247.740 60.765 248.030 60.810 ;
        RECT 248.185 60.765 248.505 60.825 ;
        RECT 247.740 60.625 248.505 60.765 ;
        RECT 247.740 60.580 248.030 60.625 ;
        RECT 248.185 60.565 248.505 60.625 ;
        RECT 254.625 60.565 254.945 60.825 ;
        RECT 255.085 60.565 255.405 60.825 ;
        RECT 255.545 60.765 255.865 60.825 ;
        RECT 258.395 60.765 258.535 61.305 ;
        RECT 269.665 61.105 269.805 61.305 ;
        RECT 279.925 61.305 283.005 61.445 ;
        RECT 279.925 61.245 280.245 61.305 ;
        RECT 282.685 61.245 283.005 61.305 ;
        RECT 284.525 61.245 284.845 61.505 ;
        RECT 285.460 61.260 285.750 61.490 ;
        RECT 287.375 61.445 287.515 61.645 ;
        RECT 287.745 61.645 288.510 61.785 ;
        RECT 287.745 61.585 288.065 61.645 ;
        RECT 288.220 61.600 288.510 61.645 ;
        RECT 288.755 61.645 300.855 61.785 ;
        RECT 301.085 61.785 301.405 61.845 ;
        RECT 308.905 61.785 309.225 61.845 ;
        RECT 301.085 61.645 309.225 61.785 ;
        RECT 288.755 61.490 288.895 61.645 ;
        RECT 301.085 61.585 301.405 61.645 ;
        RECT 308.905 61.585 309.225 61.645 ;
        RECT 288.680 61.445 288.970 61.490 ;
        RECT 287.375 61.305 288.970 61.445 ;
        RECT 288.680 61.260 288.970 61.305 ;
        RECT 280.845 61.105 281.165 61.165 ;
        RECT 269.665 60.965 281.165 61.105 ;
        RECT 280.845 60.905 281.165 60.965 ;
        RECT 281.765 61.105 282.085 61.165 ;
        RECT 285.535 61.105 285.675 61.260 ;
        RECT 289.585 61.245 289.905 61.505 ;
        RECT 297.880 61.260 298.170 61.490 ;
        RECT 298.325 61.445 298.645 61.505 ;
        RECT 301.560 61.445 301.850 61.490 ;
        RECT 298.325 61.305 301.850 61.445 ;
        RECT 289.675 61.105 289.815 61.245 ;
        RECT 281.765 60.965 289.815 61.105 ;
        RECT 296.945 61.105 297.265 61.165 ;
        RECT 297.955 61.105 298.095 61.260 ;
        RECT 298.325 61.245 298.645 61.305 ;
        RECT 301.560 61.260 301.850 61.305 ;
        RECT 302.020 61.260 302.310 61.490 ;
        RECT 302.095 61.105 302.235 61.260 ;
        RECT 296.945 60.965 302.235 61.105 ;
        RECT 281.765 60.905 282.085 60.965 ;
        RECT 296.945 60.905 297.265 60.965 ;
        RECT 255.545 60.625 258.535 60.765 ;
        RECT 260.145 60.765 260.465 60.825 ;
        RECT 260.620 60.765 260.910 60.810 ;
        RECT 260.145 60.625 260.910 60.765 ;
        RECT 255.545 60.565 255.865 60.625 ;
        RECT 260.145 60.565 260.465 60.625 ;
        RECT 260.620 60.580 260.910 60.625 ;
        RECT 284.525 60.765 284.845 60.825 ;
        RECT 286.380 60.765 286.670 60.810 ;
        RECT 284.525 60.625 286.670 60.765 ;
        RECT 284.525 60.565 284.845 60.625 ;
        RECT 286.380 60.580 286.670 60.625 ;
        RECT 299.260 60.765 299.550 60.810 ;
        RECT 302.005 60.765 302.325 60.825 ;
        RECT 299.260 60.625 302.325 60.765 ;
        RECT 299.260 60.580 299.550 60.625 ;
        RECT 302.005 60.565 302.325 60.625 ;
        RECT 162.095 59.945 311.135 60.425 ;
        RECT 221.505 59.545 221.825 59.805 ;
        RECT 239.445 59.745 239.765 59.805 ;
        RECT 239.920 59.745 240.210 59.790 ;
        RECT 239.445 59.605 240.210 59.745 ;
        RECT 239.445 59.545 239.765 59.605 ;
        RECT 239.920 59.560 240.210 59.605 ;
        RECT 252.785 59.745 253.105 59.805 ;
        RECT 259.225 59.745 259.545 59.805 ;
        RECT 261.540 59.745 261.830 59.790 ;
        RECT 252.785 59.605 261.830 59.745 ;
        RECT 252.785 59.545 253.105 59.605 ;
        RECT 259.225 59.545 259.545 59.605 ;
        RECT 261.540 59.560 261.830 59.605 ;
        RECT 287.745 59.745 288.065 59.805 ;
        RECT 301.085 59.745 301.405 59.805 ;
        RECT 287.745 59.605 292.115 59.745 ;
        RECT 287.745 59.545 288.065 59.605 ;
        RECT 176.885 59.205 177.205 59.465 ;
        RECT 179.645 59.405 179.965 59.465 ;
        RECT 177.895 59.265 179.965 59.405 ;
        RECT 177.895 58.770 178.035 59.265 ;
        RECT 179.645 59.205 179.965 59.265 ;
        RECT 181.485 59.405 181.805 59.465 ;
        RECT 184.705 59.405 185.025 59.465 ;
        RECT 187.005 59.405 187.325 59.465 ;
        RECT 188.845 59.405 189.165 59.465 ;
        RECT 191.145 59.405 191.465 59.465 ;
        RECT 181.485 59.265 185.025 59.405 ;
        RECT 181.485 59.205 181.805 59.265 ;
        RECT 184.705 59.205 185.025 59.265 ;
        RECT 185.715 59.265 189.165 59.405 ;
        RECT 178.740 59.065 179.030 59.110 ;
        RECT 183.325 59.065 183.645 59.125 ;
        RECT 185.715 59.110 185.855 59.265 ;
        RECT 187.005 59.205 187.325 59.265 ;
        RECT 188.845 59.205 189.165 59.265 ;
        RECT 189.395 59.265 191.465 59.405 ;
        RECT 178.740 58.925 183.645 59.065 ;
        RECT 178.740 58.880 179.030 58.925 ;
        RECT 177.820 58.540 178.110 58.770 ;
        RECT 172.745 58.385 173.065 58.445 ;
        RECT 178.815 58.385 178.955 58.880 ;
        RECT 183.325 58.865 183.645 58.925 ;
        RECT 183.800 59.065 184.090 59.110 ;
        RECT 183.800 58.925 185.395 59.065 ;
        RECT 183.800 58.880 184.090 58.925 ;
        RECT 181.485 58.525 181.805 58.785 ;
        RECT 184.245 58.525 184.565 58.785 ;
        RECT 185.255 58.725 185.395 58.925 ;
        RECT 185.640 58.880 185.930 59.110 ;
        RECT 188.385 59.065 188.705 59.125 ;
        RECT 189.395 59.065 189.535 59.265 ;
        RECT 191.145 59.205 191.465 59.265 ;
        RECT 196.665 59.405 196.985 59.465 ;
        RECT 197.140 59.405 197.430 59.450 ;
        RECT 196.665 59.265 197.430 59.405 ;
        RECT 196.665 59.205 196.985 59.265 ;
        RECT 197.140 59.220 197.430 59.265 ;
        RECT 201.725 59.405 202.045 59.465 ;
        RECT 203.120 59.405 203.410 59.450 ;
        RECT 201.725 59.265 203.410 59.405 ;
        RECT 201.725 59.205 202.045 59.265 ;
        RECT 203.120 59.220 203.410 59.265 ;
        RECT 213.650 59.405 213.940 59.450 ;
        RECT 215.540 59.405 215.830 59.450 ;
        RECT 218.660 59.405 218.950 59.450 ;
        RECT 213.650 59.265 218.950 59.405 ;
        RECT 213.650 59.220 213.940 59.265 ;
        RECT 215.540 59.220 215.830 59.265 ;
        RECT 218.660 59.220 218.950 59.265 ;
        RECT 232.050 59.405 232.340 59.450 ;
        RECT 233.940 59.405 234.230 59.450 ;
        RECT 237.060 59.405 237.350 59.450 ;
        RECT 232.050 59.265 237.350 59.405 ;
        RECT 232.050 59.220 232.340 59.265 ;
        RECT 233.940 59.220 234.230 59.265 ;
        RECT 237.060 59.220 237.350 59.265 ;
        RECT 245.425 59.205 245.745 59.465 ;
        RECT 291.975 59.450 292.115 59.605 ;
        RECT 297.035 59.605 301.405 59.745 ;
        RECT 253.670 59.405 253.960 59.450 ;
        RECT 255.560 59.405 255.850 59.450 ;
        RECT 258.680 59.405 258.970 59.450 ;
        RECT 253.670 59.265 258.970 59.405 ;
        RECT 253.670 59.220 253.960 59.265 ;
        RECT 255.560 59.220 255.850 59.265 ;
        RECT 258.680 59.220 258.970 59.265 ;
        RECT 284.030 59.405 284.320 59.450 ;
        RECT 285.920 59.405 286.210 59.450 ;
        RECT 289.040 59.405 289.330 59.450 ;
        RECT 284.030 59.265 289.330 59.405 ;
        RECT 284.030 59.220 284.320 59.265 ;
        RECT 285.920 59.220 286.210 59.265 ;
        RECT 289.040 59.220 289.330 59.265 ;
        RECT 291.900 59.220 292.190 59.450 ;
        RECT 293.725 59.405 294.045 59.465 ;
        RECT 297.035 59.405 297.175 59.605 ;
        RECT 301.085 59.545 301.405 59.605 ;
        RECT 293.725 59.265 297.175 59.405 ;
        RECT 297.520 59.405 297.810 59.450 ;
        RECT 300.640 59.405 300.930 59.450 ;
        RECT 302.530 59.405 302.820 59.450 ;
        RECT 297.520 59.265 302.820 59.405 ;
        RECT 293.725 59.205 294.045 59.265 ;
        RECT 297.520 59.220 297.810 59.265 ;
        RECT 300.640 59.220 300.930 59.265 ;
        RECT 302.530 59.220 302.820 59.265 ;
        RECT 188.385 58.925 189.535 59.065 ;
        RECT 188.385 58.865 188.705 58.925 ;
        RECT 190.685 58.865 191.005 59.125 ;
        RECT 193.905 58.865 194.225 59.125 ;
        RECT 195.285 58.865 195.605 59.125 ;
        RECT 202.645 58.865 202.965 59.125 ;
        RECT 210.925 59.065 211.245 59.125 ;
        RECT 203.195 58.925 211.245 59.065 ;
        RECT 186.085 58.735 186.405 58.795 ;
        RECT 185.715 58.725 186.405 58.735 ;
        RECT 185.255 58.595 186.405 58.725 ;
        RECT 185.255 58.585 185.855 58.595 ;
        RECT 186.085 58.535 186.405 58.595 ;
        RECT 186.545 58.525 186.865 58.785 ;
        RECT 187.465 58.725 187.785 58.785 ;
        RECT 187.940 58.725 188.230 58.770 ;
        RECT 191.160 58.725 191.450 58.770 ;
        RECT 187.465 58.585 188.230 58.725 ;
        RECT 187.465 58.525 187.785 58.585 ;
        RECT 187.940 58.540 188.230 58.585 ;
        RECT 188.475 58.585 191.450 58.725 ;
        RECT 172.745 58.245 178.955 58.385 ;
        RECT 184.335 58.385 184.475 58.525 ;
        RECT 188.475 58.385 188.615 58.585 ;
        RECT 191.160 58.540 191.450 58.585 ;
        RECT 191.620 58.725 191.910 58.770 ;
        RECT 192.065 58.725 192.385 58.785 ;
        RECT 191.620 58.585 192.385 58.725 ;
        RECT 191.620 58.540 191.910 58.585 ;
        RECT 192.065 58.525 192.385 58.585 ;
        RECT 192.540 58.540 192.830 58.770 ;
        RECT 184.335 58.245 188.615 58.385 ;
        RECT 190.225 58.385 190.545 58.445 ;
        RECT 192.615 58.385 192.755 58.540 ;
        RECT 190.225 58.245 192.755 58.385 ;
        RECT 195.375 58.385 195.515 58.865 ;
        RECT 195.745 58.725 196.065 58.785 ;
        RECT 196.220 58.725 196.510 58.770 ;
        RECT 195.745 58.585 196.510 58.725 ;
        RECT 195.745 58.525 196.065 58.585 ;
        RECT 196.220 58.540 196.510 58.585 ;
        RECT 199.885 58.725 200.205 58.785 ;
        RECT 202.200 58.725 202.490 58.770 ;
        RECT 203.195 58.725 203.335 58.925 ;
        RECT 210.925 58.865 211.245 58.925 ;
        RECT 212.780 59.065 213.070 59.110 ;
        RECT 214.145 59.065 214.465 59.125 ;
        RECT 212.780 58.925 214.465 59.065 ;
        RECT 212.780 58.880 213.070 58.925 ;
        RECT 214.145 58.865 214.465 58.925 ;
        RECT 220.585 59.065 220.905 59.125 ;
        RECT 224.280 59.065 224.570 59.110 ;
        RECT 220.585 58.925 224.570 59.065 ;
        RECT 220.585 58.865 220.905 58.925 ;
        RECT 224.280 58.880 224.570 58.925 ;
        RECT 225.200 59.065 225.490 59.110 ;
        RECT 225.645 59.065 225.965 59.125 ;
        RECT 225.200 58.925 225.965 59.065 ;
        RECT 225.200 58.880 225.490 58.925 ;
        RECT 225.645 58.865 225.965 58.925 ;
        RECT 232.545 58.865 232.865 59.125 ;
        RECT 242.205 59.065 242.525 59.125 ;
        RECT 248.185 59.065 248.505 59.125 ;
        RECT 242.205 58.925 248.505 59.065 ;
        RECT 242.205 58.865 242.525 58.925 ;
        RECT 248.185 58.865 248.505 58.925 ;
        RECT 252.800 59.065 253.090 59.110 ;
        RECT 254.165 59.065 254.485 59.125 ;
        RECT 252.800 58.925 254.485 59.065 ;
        RECT 252.800 58.880 253.090 58.925 ;
        RECT 254.165 58.865 254.485 58.925 ;
        RECT 257.845 59.065 258.165 59.125 ;
        RECT 262.000 59.065 262.290 59.110 ;
        RECT 257.845 58.925 262.290 59.065 ;
        RECT 257.845 58.865 258.165 58.925 ;
        RECT 262.000 58.880 262.290 58.925 ;
        RECT 264.760 59.065 265.050 59.110 ;
        RECT 270.740 59.065 271.030 59.110 ;
        RECT 264.760 58.925 271.030 59.065 ;
        RECT 264.760 58.880 265.050 58.925 ;
        RECT 270.740 58.880 271.030 58.925 ;
        RECT 271.200 59.065 271.490 59.110 ;
        RECT 279.925 59.065 280.245 59.125 ;
        RECT 271.200 58.925 280.245 59.065 ;
        RECT 271.200 58.880 271.490 58.925 ;
        RECT 199.885 58.585 203.335 58.725 ;
        RECT 199.885 58.525 200.205 58.585 ;
        RECT 202.200 58.540 202.490 58.585 ;
        RECT 203.565 58.525 203.885 58.785 ;
        RECT 213.245 58.725 213.535 58.770 ;
        RECT 215.080 58.725 215.370 58.770 ;
        RECT 218.660 58.725 218.950 58.770 ;
        RECT 213.245 58.585 218.950 58.725 ;
        RECT 213.245 58.540 213.535 58.585 ;
        RECT 215.080 58.540 215.370 58.585 ;
        RECT 218.660 58.540 218.950 58.585 ;
        RECT 210.005 58.385 210.325 58.445 ;
        RECT 219.740 58.430 220.030 58.745 ;
        RECT 227.485 58.525 227.805 58.785 ;
        RECT 227.945 58.725 228.265 58.785 ;
        RECT 231.180 58.725 231.470 58.770 ;
        RECT 227.945 58.585 231.470 58.725 ;
        RECT 227.945 58.525 228.265 58.585 ;
        RECT 231.180 58.540 231.470 58.585 ;
        RECT 231.645 58.725 231.935 58.770 ;
        RECT 233.480 58.725 233.770 58.770 ;
        RECT 237.060 58.725 237.350 58.770 ;
        RECT 231.645 58.585 237.350 58.725 ;
        RECT 231.645 58.540 231.935 58.585 ;
        RECT 233.480 58.540 233.770 58.585 ;
        RECT 237.060 58.540 237.350 58.585 ;
        RECT 195.375 58.245 210.325 58.385 ;
        RECT 172.745 58.185 173.065 58.245 ;
        RECT 190.225 58.185 190.545 58.245 ;
        RECT 210.005 58.185 210.325 58.245 ;
        RECT 214.160 58.200 214.450 58.430 ;
        RECT 216.440 58.385 217.090 58.430 ;
        RECT 219.740 58.385 220.330 58.430 ;
        RECT 222.885 58.385 223.205 58.445 ;
        RECT 216.440 58.245 223.205 58.385 ;
        RECT 216.440 58.200 217.090 58.245 ;
        RECT 220.040 58.200 220.330 58.245 ;
        RECT 182.420 58.045 182.710 58.090 ;
        RECT 182.865 58.045 183.185 58.105 ;
        RECT 182.420 57.905 183.185 58.045 ;
        RECT 182.420 57.860 182.710 57.905 ;
        RECT 182.865 57.845 183.185 57.905 ;
        RECT 184.705 58.045 185.025 58.105 ;
        RECT 188.845 58.045 189.165 58.105 ;
        RECT 190.315 58.045 190.455 58.185 ;
        RECT 184.705 57.905 190.455 58.045 ;
        RECT 201.280 58.045 201.570 58.090 ;
        RECT 201.725 58.045 202.045 58.105 ;
        RECT 201.280 57.905 202.045 58.045 ;
        RECT 214.235 58.045 214.375 58.200 ;
        RECT 222.885 58.185 223.205 58.245 ;
        RECT 223.820 58.385 224.110 58.430 ;
        RECT 224.725 58.385 225.045 58.445 ;
        RECT 223.820 58.245 225.045 58.385 ;
        RECT 223.820 58.200 224.110 58.245 ;
        RECT 224.725 58.185 225.045 58.245 ;
        RECT 229.325 58.385 229.645 58.445 ;
        RECT 238.140 58.430 238.430 58.745 ;
        RECT 243.600 58.725 243.890 58.770 ;
        RECT 246.345 58.725 246.665 58.785 ;
        RECT 243.600 58.585 246.665 58.725 ;
        RECT 243.600 58.540 243.890 58.585 ;
        RECT 246.345 58.525 246.665 58.585 ;
        RECT 253.265 58.725 253.555 58.770 ;
        RECT 255.100 58.725 255.390 58.770 ;
        RECT 258.680 58.725 258.970 58.770 ;
        RECT 253.265 58.585 258.970 58.725 ;
        RECT 253.265 58.540 253.555 58.585 ;
        RECT 255.100 58.540 255.390 58.585 ;
        RECT 258.680 58.540 258.970 58.585 ;
        RECT 234.840 58.385 235.490 58.430 ;
        RECT 238.140 58.385 238.730 58.430 ;
        RECT 229.325 58.245 238.730 58.385 ;
        RECT 229.325 58.185 229.645 58.245 ;
        RECT 234.840 58.200 235.490 58.245 ;
        RECT 238.440 58.200 238.730 58.245 ;
        RECT 242.665 58.385 242.985 58.445 ;
        RECT 244.645 58.385 244.935 58.430 ;
        RECT 245.885 58.385 246.205 58.445 ;
        RECT 242.665 58.245 246.205 58.385 ;
        RECT 242.665 58.185 242.985 58.245 ;
        RECT 244.645 58.200 244.935 58.245 ;
        RECT 245.885 58.185 246.205 58.245 ;
        RECT 254.180 58.385 254.470 58.430 ;
        RECT 254.625 58.385 254.945 58.445 ;
        RECT 259.760 58.430 260.050 58.745 ;
        RECT 262.905 58.525 263.225 58.785 ;
        RECT 263.365 58.525 263.685 58.785 ;
        RECT 254.180 58.245 254.945 58.385 ;
        RECT 254.180 58.200 254.470 58.245 ;
        RECT 254.625 58.185 254.945 58.245 ;
        RECT 256.460 58.385 257.110 58.430 ;
        RECT 259.760 58.385 260.350 58.430 ;
        RECT 260.605 58.385 260.925 58.445 ;
        RECT 264.835 58.385 264.975 58.880 ;
        RECT 279.925 58.865 280.245 58.925 ;
        RECT 280.845 58.865 281.165 59.125 ;
        RECT 281.765 58.865 282.085 59.125 ;
        RECT 283.160 59.065 283.450 59.110 ;
        RECT 290.505 59.065 290.825 59.125 ;
        RECT 303.400 59.065 303.690 59.110 ;
        RECT 308.905 59.065 309.225 59.125 ;
        RECT 283.160 58.925 309.225 59.065 ;
        RECT 283.160 58.880 283.450 58.925 ;
        RECT 290.505 58.865 290.825 58.925 ;
        RECT 303.400 58.880 303.690 58.925 ;
        RECT 308.905 58.865 309.225 58.925 ;
        RECT 273.040 58.725 273.330 58.770 ;
        RECT 274.405 58.725 274.725 58.785 ;
        RECT 273.040 58.585 274.725 58.725 ;
        RECT 273.040 58.540 273.330 58.585 ;
        RECT 274.405 58.525 274.725 58.585 ;
        RECT 276.245 58.725 276.565 58.785 ;
        RECT 280.400 58.725 280.690 58.770 ;
        RECT 282.685 58.725 283.005 58.785 ;
        RECT 276.245 58.585 280.155 58.725 ;
        RECT 276.245 58.525 276.565 58.585 ;
        RECT 256.460 58.245 260.925 58.385 ;
        RECT 256.460 58.200 257.110 58.245 ;
        RECT 260.060 58.200 260.350 58.245 ;
        RECT 260.605 58.185 260.925 58.245 ;
        RECT 261.155 58.245 264.975 58.385 ;
        RECT 218.285 58.045 218.605 58.105 ;
        RECT 214.235 57.905 218.605 58.045 ;
        RECT 184.705 57.845 185.025 57.905 ;
        RECT 188.845 57.845 189.165 57.905 ;
        RECT 201.280 57.860 201.570 57.905 ;
        RECT 201.725 57.845 202.045 57.905 ;
        RECT 218.285 57.845 218.605 57.905 ;
        RECT 221.980 58.045 222.270 58.090 ;
        RECT 222.425 58.045 222.745 58.105 ;
        RECT 221.980 57.905 222.745 58.045 ;
        RECT 221.980 57.860 222.270 57.905 ;
        RECT 222.425 57.845 222.745 57.905 ;
        RECT 230.720 58.045 231.010 58.090 ;
        RECT 239.445 58.045 239.765 58.105 ;
        RECT 230.720 57.905 239.765 58.045 ;
        RECT 230.720 57.860 231.010 57.905 ;
        RECT 239.445 57.845 239.765 57.905 ;
        RECT 243.585 58.045 243.905 58.105 ;
        RECT 244.060 58.045 244.350 58.090 ;
        RECT 243.585 57.905 244.350 58.045 ;
        RECT 243.585 57.845 243.905 57.905 ;
        RECT 244.060 57.860 244.350 57.905 ;
        RECT 248.185 58.045 248.505 58.105 ;
        RECT 261.155 58.045 261.295 58.245 ;
        RECT 273.500 58.200 273.790 58.430 ;
        RECT 248.185 57.905 261.295 58.045 ;
        RECT 263.840 58.045 264.130 58.090 ;
        RECT 264.285 58.045 264.605 58.105 ;
        RECT 273.575 58.045 273.715 58.200 ;
        RECT 263.840 57.905 273.715 58.045 ;
        RECT 276.705 58.045 277.025 58.105 ;
        RECT 278.560 58.045 278.850 58.090 ;
        RECT 276.705 57.905 278.850 58.045 ;
        RECT 280.015 58.045 280.155 58.585 ;
        RECT 280.400 58.585 283.005 58.725 ;
        RECT 280.400 58.540 280.690 58.585 ;
        RECT 282.685 58.525 283.005 58.585 ;
        RECT 283.625 58.725 283.915 58.770 ;
        RECT 285.460 58.725 285.750 58.770 ;
        RECT 289.040 58.725 289.330 58.770 ;
        RECT 283.625 58.585 289.330 58.725 ;
        RECT 283.625 58.540 283.915 58.585 ;
        RECT 285.460 58.540 285.750 58.585 ;
        RECT 289.040 58.540 289.330 58.585 ;
        RECT 280.845 58.385 281.165 58.445 ;
        RECT 280.845 58.245 284.295 58.385 ;
        RECT 280.845 58.185 281.165 58.245 ;
        RECT 283.605 58.045 283.925 58.105 ;
        RECT 280.015 57.905 283.925 58.045 ;
        RECT 284.155 58.045 284.295 58.245 ;
        RECT 284.525 58.185 284.845 58.445 ;
        RECT 286.825 58.430 287.145 58.445 ;
        RECT 290.120 58.430 290.410 58.745 ;
        RECT 296.440 58.430 296.730 58.745 ;
        RECT 297.520 58.725 297.810 58.770 ;
        RECT 301.100 58.725 301.390 58.770 ;
        RECT 302.935 58.725 303.225 58.770 ;
        RECT 297.520 58.585 303.225 58.725 ;
        RECT 297.520 58.540 297.810 58.585 ;
        RECT 301.100 58.540 301.390 58.585 ;
        RECT 302.935 58.540 303.225 58.585 ;
        RECT 286.820 58.385 287.470 58.430 ;
        RECT 290.120 58.385 290.710 58.430 ;
        RECT 296.140 58.385 296.730 58.430 ;
        RECT 299.380 58.385 300.030 58.430 ;
        RECT 286.455 58.245 290.710 58.385 ;
        RECT 286.455 58.045 286.595 58.245 ;
        RECT 286.820 58.200 287.470 58.245 ;
        RECT 290.420 58.200 290.710 58.245 ;
        RECT 291.055 58.245 300.030 58.385 ;
        RECT 286.825 58.185 287.145 58.200 ;
        RECT 291.055 58.045 291.195 58.245 ;
        RECT 284.155 57.905 291.195 58.045 ;
        RECT 293.725 58.045 294.045 58.105 ;
        RECT 294.660 58.045 294.950 58.090 ;
        RECT 293.725 57.905 294.950 58.045 ;
        RECT 295.655 58.045 295.795 58.245 ;
        RECT 296.140 58.200 296.430 58.245 ;
        RECT 299.380 58.200 300.030 58.245 ;
        RECT 302.005 58.185 302.325 58.445 ;
        RECT 297.865 58.045 298.185 58.105 ;
        RECT 295.655 57.905 298.185 58.045 ;
        RECT 248.185 57.845 248.505 57.905 ;
        RECT 263.840 57.860 264.130 57.905 ;
        RECT 264.285 57.845 264.605 57.905 ;
        RECT 276.705 57.845 277.025 57.905 ;
        RECT 278.560 57.860 278.850 57.905 ;
        RECT 283.605 57.845 283.925 57.905 ;
        RECT 293.725 57.845 294.045 57.905 ;
        RECT 294.660 57.860 294.950 57.905 ;
        RECT 297.865 57.845 298.185 57.905 ;
        RECT 162.095 57.225 311.135 57.705 ;
        RECT 164.925 57.025 165.245 57.085 ;
        RECT 172.300 57.025 172.590 57.070 ;
        RECT 175.060 57.025 175.350 57.070 ;
        RECT 175.965 57.025 176.285 57.085 ;
        RECT 164.925 56.885 176.285 57.025 ;
        RECT 164.925 56.825 165.245 56.885 ;
        RECT 172.300 56.840 172.590 56.885 ;
        RECT 175.060 56.840 175.350 56.885 ;
        RECT 175.965 56.825 176.285 56.885 ;
        RECT 184.245 56.825 184.565 57.085 ;
        RECT 186.545 57.025 186.865 57.085 ;
        RECT 187.925 57.025 188.245 57.085 ;
        RECT 186.545 56.885 188.245 57.025 ;
        RECT 186.545 56.825 186.865 56.885 ;
        RECT 187.925 56.825 188.245 56.885 ;
        RECT 189.765 57.025 190.085 57.085 ;
        RECT 192.080 57.025 192.370 57.070 ;
        RECT 189.765 56.885 192.370 57.025 ;
        RECT 189.765 56.825 190.085 56.885 ;
        RECT 192.080 56.840 192.370 56.885 ;
        RECT 203.105 57.025 203.425 57.085 ;
        RECT 203.580 57.025 203.870 57.070 ;
        RECT 203.105 56.885 203.870 57.025 ;
        RECT 203.105 56.825 203.425 56.885 ;
        RECT 203.580 56.840 203.870 56.885 ;
        RECT 208.625 57.025 208.945 57.085 ;
        RECT 209.100 57.025 209.390 57.070 ;
        RECT 213.240 57.025 213.530 57.070 ;
        RECT 215.525 57.025 215.845 57.085 ;
        RECT 208.625 56.885 209.390 57.025 ;
        RECT 208.625 56.825 208.945 56.885 ;
        RECT 209.100 56.840 209.390 56.885 ;
        RECT 211.475 56.885 212.995 57.025 ;
        RECT 172.745 56.485 173.065 56.745 ;
        RECT 174.585 56.685 174.905 56.745 ;
        RECT 179.660 56.685 179.950 56.730 ;
        RECT 174.585 56.545 179.950 56.685 ;
        RECT 174.585 56.485 174.905 56.545 ;
        RECT 179.660 56.500 179.950 56.545 ;
        RECT 189.195 56.500 189.485 56.730 ;
        RECT 195.760 56.685 196.050 56.730 ;
        RECT 196.205 56.685 196.525 56.745 ;
        RECT 198.045 56.730 198.365 56.745 ;
        RECT 195.760 56.545 196.525 56.685 ;
        RECT 195.760 56.500 196.050 56.545 ;
        RECT 175.965 56.145 176.285 56.405 ;
        RECT 176.425 56.345 176.745 56.405 ;
        RECT 176.900 56.345 177.190 56.390 ;
        RECT 176.425 56.205 177.190 56.345 ;
        RECT 176.425 56.145 176.745 56.205 ;
        RECT 176.900 56.160 177.190 56.205 ;
        RECT 177.820 56.345 178.110 56.390 ;
        RECT 179.185 56.345 179.505 56.405 ;
        RECT 177.820 56.205 179.505 56.345 ;
        RECT 177.820 56.160 178.110 56.205 ;
        RECT 179.185 56.145 179.505 56.205 ;
        RECT 180.565 56.345 180.885 56.405 ;
        RECT 181.500 56.345 181.790 56.390 ;
        RECT 185.165 56.345 185.485 56.405 ;
        RECT 180.565 56.205 185.485 56.345 ;
        RECT 180.565 56.145 180.885 56.205 ;
        RECT 181.500 56.160 181.790 56.205 ;
        RECT 185.165 56.145 185.485 56.205 ;
        RECT 185.635 56.160 185.925 56.390 ;
        RECT 173.665 55.805 173.985 56.065 ;
        RECT 175.505 56.005 175.825 56.065 ;
        RECT 178.740 56.005 179.030 56.050 ;
        RECT 175.505 55.865 179.030 56.005 ;
        RECT 175.505 55.805 175.825 55.865 ;
        RECT 178.740 55.820 179.030 55.865 ;
        RECT 184.705 55.665 185.025 55.725 ;
        RECT 185.715 55.665 185.855 56.160 ;
        RECT 186.085 56.145 186.405 56.405 ;
        RECT 189.270 56.345 189.410 56.500 ;
        RECT 196.205 56.485 196.525 56.545 ;
        RECT 198.040 56.685 198.690 56.730 ;
        RECT 201.640 56.685 201.930 56.730 ;
        RECT 198.040 56.545 201.930 56.685 ;
        RECT 198.040 56.500 198.690 56.545 ;
        RECT 201.340 56.500 201.930 56.545 ;
        RECT 205.420 56.685 205.710 56.730 ;
        RECT 206.785 56.685 207.105 56.745 ;
        RECT 211.475 56.730 211.615 56.885 ;
        RECT 210.940 56.685 211.230 56.730 ;
        RECT 211.400 56.685 211.690 56.730 ;
        RECT 205.420 56.545 211.690 56.685 ;
        RECT 205.420 56.500 205.710 56.545 ;
        RECT 198.045 56.485 198.365 56.500 ;
        RECT 188.935 56.205 189.410 56.345 ;
        RECT 191.145 56.345 191.465 56.405 ;
        RECT 193.000 56.345 193.290 56.390 ;
        RECT 191.145 56.205 193.290 56.345 ;
        RECT 188.935 56.065 189.075 56.205 ;
        RECT 191.145 56.145 191.465 56.205 ;
        RECT 193.000 56.160 193.290 56.205 ;
        RECT 194.845 56.345 195.135 56.390 ;
        RECT 196.680 56.345 196.970 56.390 ;
        RECT 200.260 56.345 200.550 56.390 ;
        RECT 194.845 56.205 200.550 56.345 ;
        RECT 194.845 56.160 195.135 56.205 ;
        RECT 196.680 56.160 196.970 56.205 ;
        RECT 200.260 56.160 200.550 56.205 ;
        RECT 201.340 56.185 201.630 56.500 ;
        RECT 206.785 56.485 207.105 56.545 ;
        RECT 210.940 56.500 211.230 56.545 ;
        RECT 211.400 56.500 211.690 56.545 ;
        RECT 212.320 56.500 212.610 56.730 ;
        RECT 212.855 56.685 212.995 56.885 ;
        RECT 213.240 56.885 215.845 57.025 ;
        RECT 213.240 56.840 213.530 56.885 ;
        RECT 215.525 56.825 215.845 56.885 ;
        RECT 218.300 57.025 218.590 57.070 ;
        RECT 218.745 57.025 219.065 57.085 ;
        RECT 263.840 57.025 264.130 57.070 ;
        RECT 267.965 57.025 268.285 57.085 ;
        RECT 218.300 56.885 247.495 57.025 ;
        RECT 218.300 56.840 218.590 56.885 ;
        RECT 218.745 56.825 219.065 56.885 ;
        RECT 219.205 56.685 219.525 56.745 ;
        RECT 222.885 56.730 223.205 56.745 ;
        RECT 212.855 56.545 219.525 56.685 ;
        RECT 204.485 56.345 204.805 56.405 ;
        RECT 203.195 56.205 204.805 56.345 ;
        RECT 188.845 55.805 189.165 56.065 ;
        RECT 189.780 55.820 190.070 56.050 ;
        RECT 190.240 56.005 190.530 56.050 ;
        RECT 190.685 56.005 191.005 56.065 ;
        RECT 190.240 55.865 191.005 56.005 ;
        RECT 190.240 55.820 190.530 55.865 ;
        RECT 189.855 55.665 189.995 55.820 ;
        RECT 190.685 55.805 191.005 55.865 ;
        RECT 191.620 56.005 191.910 56.050 ;
        RECT 192.065 56.005 192.385 56.065 ;
        RECT 191.620 55.865 192.385 56.005 ;
        RECT 191.620 55.820 191.910 55.865 ;
        RECT 192.065 55.805 192.385 55.865 ;
        RECT 193.905 56.005 194.225 56.065 ;
        RECT 203.195 56.050 203.335 56.205 ;
        RECT 204.485 56.145 204.805 56.205 ;
        RECT 209.545 56.345 209.865 56.405 ;
        RECT 210.020 56.345 210.310 56.390 ;
        RECT 209.545 56.205 210.310 56.345 ;
        RECT 212.395 56.345 212.535 56.500 ;
        RECT 219.205 56.485 219.525 56.545 ;
        RECT 219.780 56.685 220.070 56.730 ;
        RECT 222.885 56.685 223.670 56.730 ;
        RECT 219.780 56.545 223.670 56.685 ;
        RECT 219.780 56.500 220.370 56.545 ;
        RECT 213.225 56.345 213.545 56.405 ;
        RECT 212.395 56.205 213.545 56.345 ;
        RECT 209.545 56.145 209.865 56.205 ;
        RECT 210.020 56.160 210.310 56.205 ;
        RECT 213.225 56.145 213.545 56.205 ;
        RECT 215.030 56.160 215.320 56.390 ;
        RECT 194.380 56.005 194.670 56.050 ;
        RECT 193.905 55.865 194.670 56.005 ;
        RECT 193.905 55.805 194.225 55.865 ;
        RECT 194.380 55.820 194.670 55.865 ;
        RECT 203.120 55.820 203.410 56.050 ;
        RECT 184.705 55.525 189.995 55.665 ;
        RECT 195.250 55.665 195.540 55.710 ;
        RECT 197.140 55.665 197.430 55.710 ;
        RECT 200.260 55.665 200.550 55.710 ;
        RECT 195.250 55.525 200.550 55.665 ;
        RECT 184.705 55.465 185.025 55.525 ;
        RECT 195.250 55.480 195.540 55.525 ;
        RECT 197.140 55.480 197.430 55.525 ;
        RECT 200.260 55.480 200.550 55.525 ;
        RECT 210.925 55.665 211.245 55.725 ;
        RECT 215.105 55.665 215.245 56.160 ;
        RECT 215.985 56.145 216.305 56.405 ;
        RECT 216.460 56.345 216.750 56.390 ;
        RECT 218.285 56.345 218.605 56.405 ;
        RECT 216.460 56.205 218.605 56.345 ;
        RECT 216.460 56.160 216.750 56.205 ;
        RECT 218.285 56.145 218.605 56.205 ;
        RECT 220.080 56.185 220.370 56.500 ;
        RECT 222.885 56.500 223.670 56.545 ;
        RECT 225.185 56.685 225.505 56.745 ;
        RECT 225.660 56.685 225.950 56.730 ;
        RECT 225.185 56.545 225.950 56.685 ;
        RECT 222.885 56.485 223.205 56.500 ;
        RECT 225.185 56.485 225.505 56.545 ;
        RECT 225.660 56.500 225.950 56.545 ;
        RECT 228.865 56.485 229.185 56.745 ;
        RECT 229.325 56.685 229.645 56.745 ;
        RECT 231.160 56.685 231.810 56.730 ;
        RECT 234.760 56.685 235.050 56.730 ;
        RECT 245.440 56.685 245.730 56.730 ;
        RECT 229.325 56.545 235.050 56.685 ;
        RECT 229.325 56.485 229.645 56.545 ;
        RECT 231.160 56.500 231.810 56.545 ;
        RECT 234.460 56.500 235.050 56.545 ;
        RECT 236.775 56.545 245.730 56.685 ;
        RECT 221.160 56.345 221.450 56.390 ;
        RECT 224.740 56.345 225.030 56.390 ;
        RECT 226.575 56.345 226.865 56.390 ;
        RECT 221.160 56.205 226.865 56.345 ;
        RECT 221.160 56.160 221.450 56.205 ;
        RECT 224.740 56.160 225.030 56.205 ;
        RECT 226.575 56.160 226.865 56.205 ;
        RECT 227.040 56.345 227.330 56.390 ;
        RECT 227.485 56.345 227.805 56.405 ;
        RECT 227.040 56.205 227.805 56.345 ;
        RECT 227.040 56.160 227.330 56.205 ;
        RECT 227.485 56.145 227.805 56.205 ;
        RECT 227.965 56.345 228.255 56.390 ;
        RECT 229.800 56.345 230.090 56.390 ;
        RECT 233.380 56.345 233.670 56.390 ;
        RECT 227.965 56.205 233.670 56.345 ;
        RECT 227.965 56.160 228.255 56.205 ;
        RECT 229.800 56.160 230.090 56.205 ;
        RECT 233.380 56.160 233.670 56.205 ;
        RECT 234.460 56.185 234.750 56.500 ;
        RECT 236.775 56.390 236.915 56.545 ;
        RECT 245.440 56.500 245.730 56.545 ;
        RECT 236.700 56.160 236.990 56.390 ;
        RECT 237.620 56.345 237.910 56.390 ;
        RECT 238.985 56.345 239.305 56.405 ;
        RECT 237.620 56.205 239.305 56.345 ;
        RECT 237.620 56.160 237.910 56.205 ;
        RECT 215.540 56.005 215.830 56.050 ;
        RECT 216.075 56.005 216.215 56.145 ;
        RECT 215.540 55.865 216.215 56.005 ;
        RECT 230.705 56.005 231.025 56.065 ;
        RECT 236.240 56.005 236.530 56.050 ;
        RECT 230.705 55.865 236.530 56.005 ;
        RECT 215.540 55.820 215.830 55.865 ;
        RECT 230.705 55.805 231.025 55.865 ;
        RECT 236.240 55.820 236.530 55.865 ;
        RECT 210.925 55.525 215.245 55.665 ;
        RECT 210.925 55.465 211.245 55.525 ;
        RECT 215.985 55.465 216.305 55.725 ;
        RECT 221.160 55.665 221.450 55.710 ;
        RECT 224.280 55.665 224.570 55.710 ;
        RECT 226.170 55.665 226.460 55.710 ;
        RECT 221.160 55.525 226.460 55.665 ;
        RECT 221.160 55.480 221.450 55.525 ;
        RECT 224.280 55.480 224.570 55.525 ;
        RECT 226.170 55.480 226.460 55.525 ;
        RECT 228.370 55.665 228.660 55.710 ;
        RECT 230.260 55.665 230.550 55.710 ;
        RECT 233.380 55.665 233.670 55.710 ;
        RECT 236.775 55.665 236.915 56.160 ;
        RECT 238.985 56.145 239.305 56.205 ;
        RECT 242.205 56.345 242.525 56.405 ;
        RECT 244.520 56.345 244.810 56.390 ;
        RECT 242.205 56.205 244.810 56.345 ;
        RECT 242.205 56.145 242.525 56.205 ;
        RECT 244.520 56.160 244.810 56.205 ;
        RECT 238.065 56.005 238.385 56.065 ;
        RECT 242.680 56.005 242.970 56.050 ;
        RECT 238.065 55.865 242.970 56.005 ;
        RECT 245.515 56.005 245.655 56.500 ;
        RECT 247.355 56.390 247.495 56.885 ;
        RECT 253.795 56.885 268.285 57.025 ;
        RECT 248.185 56.685 248.505 56.745 ;
        RECT 252.785 56.685 253.105 56.745 ;
        RECT 248.185 56.545 253.105 56.685 ;
        RECT 248.185 56.485 248.505 56.545 ;
        RECT 252.785 56.485 253.105 56.545 ;
        RECT 247.280 56.160 247.570 56.390 ;
        RECT 247.725 56.345 248.045 56.405 ;
        RECT 251.880 56.345 252.170 56.390 ;
        RECT 247.725 56.205 252.170 56.345 ;
        RECT 247.725 56.145 248.045 56.205 ;
        RECT 251.880 56.160 252.170 56.205 ;
        RECT 252.325 56.145 252.645 56.405 ;
        RECT 253.795 56.390 253.935 56.885 ;
        RECT 263.840 56.840 264.130 56.885 ;
        RECT 267.965 56.825 268.285 56.885 ;
        RECT 278.545 57.025 278.865 57.085 ;
        RECT 278.545 56.885 283.375 57.025 ;
        RECT 278.545 56.825 278.865 56.885 ;
        RECT 255.085 56.685 255.405 56.745 ;
        RECT 255.560 56.685 255.850 56.730 ;
        RECT 255.085 56.545 255.850 56.685 ;
        RECT 255.085 56.485 255.405 56.545 ;
        RECT 255.560 56.500 255.850 56.545 ;
        RECT 257.840 56.685 258.490 56.730 ;
        RECT 260.605 56.685 260.925 56.745 ;
        RECT 261.440 56.685 261.730 56.730 ;
        RECT 257.840 56.545 261.730 56.685 ;
        RECT 257.840 56.500 258.490 56.545 ;
        RECT 260.605 56.485 260.925 56.545 ;
        RECT 261.140 56.500 261.730 56.545 ;
        RECT 262.905 56.685 263.225 56.745 ;
        RECT 276.245 56.685 276.565 56.745 ;
        RECT 262.905 56.545 276.565 56.685 ;
        RECT 253.720 56.160 254.010 56.390 ;
        RECT 254.645 56.345 254.935 56.390 ;
        RECT 256.480 56.345 256.770 56.390 ;
        RECT 260.060 56.345 260.350 56.390 ;
        RECT 254.645 56.205 260.350 56.345 ;
        RECT 254.645 56.160 254.935 56.205 ;
        RECT 256.480 56.160 256.770 56.205 ;
        RECT 260.060 56.160 260.350 56.205 ;
        RECT 261.140 56.185 261.430 56.500 ;
        RECT 262.905 56.485 263.225 56.545 ;
        RECT 276.245 56.485 276.565 56.545 ;
        RECT 276.705 56.485 277.025 56.745 ;
        RECT 278.085 56.685 278.405 56.745 ;
        RECT 279.005 56.730 279.325 56.745 ;
        RECT 279.000 56.685 279.650 56.730 ;
        RECT 282.600 56.685 282.890 56.730 ;
        RECT 278.085 56.545 282.890 56.685 ;
        RECT 283.235 56.685 283.375 56.885 ;
        RECT 284.065 56.825 284.385 57.085 ;
        RECT 292.805 57.025 293.125 57.085 ;
        RECT 293.280 57.025 293.570 57.070 ;
        RECT 284.615 56.885 293.570 57.025 ;
        RECT 284.615 56.685 284.755 56.885 ;
        RECT 292.805 56.825 293.125 56.885 ;
        RECT 293.280 56.840 293.570 56.885 ;
        RECT 293.740 57.025 294.030 57.070 ;
        RECT 296.025 57.025 296.345 57.085 ;
        RECT 293.740 56.885 296.345 57.025 ;
        RECT 293.740 56.840 294.030 56.885 ;
        RECT 296.025 56.825 296.345 56.885 ;
        RECT 283.235 56.545 284.755 56.685 ;
        RECT 288.205 56.685 288.525 56.745 ;
        RECT 289.140 56.685 289.430 56.730 ;
        RECT 288.205 56.545 289.430 56.685 ;
        RECT 278.085 56.485 278.405 56.545 ;
        RECT 279.000 56.500 279.650 56.545 ;
        RECT 282.300 56.500 282.890 56.545 ;
        RECT 279.005 56.485 279.325 56.500 ;
        RECT 263.380 56.345 263.670 56.390 ;
        RECT 264.745 56.345 265.065 56.405 ;
        RECT 263.380 56.205 265.065 56.345 ;
        RECT 263.380 56.160 263.670 56.205 ;
        RECT 264.745 56.145 265.065 56.205 ;
        RECT 275.805 56.345 276.095 56.390 ;
        RECT 277.640 56.345 277.930 56.390 ;
        RECT 281.220 56.345 281.510 56.390 ;
        RECT 275.805 56.205 281.510 56.345 ;
        RECT 275.805 56.160 276.095 56.205 ;
        RECT 277.640 56.160 277.930 56.205 ;
        RECT 281.220 56.160 281.510 56.205 ;
        RECT 282.300 56.185 282.590 56.500 ;
        RECT 288.205 56.485 288.525 56.545 ;
        RECT 289.140 56.500 289.430 56.545 ;
        RECT 289.585 56.685 289.905 56.745 ;
        RECT 297.865 56.685 298.185 56.745 ;
        RECT 302.020 56.685 302.310 56.730 ;
        RECT 305.240 56.685 305.530 56.730 ;
        RECT 289.585 56.545 294.415 56.685 ;
        RECT 289.585 56.485 289.905 56.545 ;
        RECT 283.605 56.345 283.925 56.405 ;
        RECT 293.725 56.345 294.045 56.405 ;
        RECT 283.605 56.205 294.045 56.345 ;
        RECT 283.605 56.145 283.925 56.205 ;
        RECT 293.725 56.145 294.045 56.205 ;
        RECT 250.945 56.005 251.265 56.065 ;
        RECT 245.515 55.865 251.265 56.005 ;
        RECT 238.065 55.805 238.385 55.865 ;
        RECT 242.680 55.820 242.970 55.865 ;
        RECT 250.945 55.805 251.265 55.865 ;
        RECT 254.165 55.805 254.485 56.065 ;
        RECT 257.845 56.005 258.165 56.065 ;
        RECT 254.715 55.865 258.165 56.005 ;
        RECT 228.370 55.525 233.670 55.665 ;
        RECT 228.370 55.480 228.660 55.525 ;
        RECT 230.260 55.480 230.550 55.525 ;
        RECT 233.380 55.480 233.670 55.525 ;
        RECT 236.315 55.525 236.915 55.665 ;
        RECT 238.540 55.665 238.830 55.710 ;
        RECT 243.125 55.665 243.445 55.725 ;
        RECT 238.540 55.525 243.445 55.665 ;
        RECT 167.225 55.325 167.545 55.385 ;
        RECT 170.460 55.325 170.750 55.370 ;
        RECT 167.225 55.185 170.750 55.325 ;
        RECT 167.225 55.125 167.545 55.185 ;
        RECT 170.460 55.140 170.750 55.185 ;
        RECT 179.645 55.325 179.965 55.385 ;
        RECT 187.925 55.325 188.245 55.385 ;
        RECT 188.400 55.325 188.690 55.370 ;
        RECT 195.745 55.325 196.065 55.385 ;
        RECT 179.645 55.185 196.065 55.325 ;
        RECT 179.645 55.125 179.965 55.185 ;
        RECT 187.925 55.125 188.245 55.185 ;
        RECT 188.400 55.140 188.690 55.185 ;
        RECT 195.745 55.125 196.065 55.185 ;
        RECT 214.160 55.325 214.450 55.370 ;
        RECT 215.065 55.325 215.385 55.385 ;
        RECT 214.160 55.185 215.385 55.325 ;
        RECT 214.160 55.140 214.450 55.185 ;
        RECT 215.065 55.125 215.385 55.185 ;
        RECT 223.805 55.325 224.125 55.385 ;
        RECT 236.315 55.325 236.455 55.525 ;
        RECT 238.540 55.480 238.830 55.525 ;
        RECT 243.125 55.465 243.445 55.525 ;
        RECT 250.500 55.665 250.790 55.710 ;
        RECT 254.715 55.665 254.855 55.865 ;
        RECT 257.845 55.805 258.165 55.865 ;
        RECT 275.325 55.805 275.645 56.065 ;
        RECT 284.065 56.005 284.385 56.065 ;
        RECT 275.875 55.865 284.385 56.005 ;
        RECT 250.500 55.525 254.855 55.665 ;
        RECT 255.050 55.665 255.340 55.710 ;
        RECT 256.940 55.665 257.230 55.710 ;
        RECT 260.060 55.665 260.350 55.710 ;
        RECT 255.050 55.525 260.350 55.665 ;
        RECT 250.500 55.480 250.790 55.525 ;
        RECT 255.050 55.480 255.340 55.525 ;
        RECT 256.940 55.480 257.230 55.525 ;
        RECT 260.060 55.480 260.350 55.525 ;
        RECT 262.445 55.665 262.765 55.725 ;
        RECT 262.920 55.665 263.210 55.710 ;
        RECT 262.445 55.525 263.210 55.665 ;
        RECT 262.445 55.465 262.765 55.525 ;
        RECT 262.920 55.480 263.210 55.525 ;
        RECT 263.365 55.665 263.685 55.725 ;
        RECT 275.875 55.665 276.015 55.865 ;
        RECT 284.065 55.805 284.385 55.865 ;
        RECT 285.460 56.005 285.750 56.050 ;
        RECT 285.905 56.005 286.225 56.065 ;
        RECT 294.275 56.050 294.415 56.545 ;
        RECT 297.865 56.545 305.530 56.685 ;
        RECT 297.865 56.485 298.185 56.545 ;
        RECT 302.020 56.500 302.310 56.545 ;
        RECT 305.240 56.500 305.530 56.545 ;
        RECT 306.160 56.685 306.450 56.730 ;
        RECT 308.000 56.685 308.290 56.730 ;
        RECT 306.160 56.545 308.290 56.685 ;
        RECT 306.160 56.500 306.450 56.545 ;
        RECT 308.000 56.500 308.290 56.545 ;
        RECT 303.840 56.345 304.130 56.390 ;
        RECT 306.160 56.345 306.375 56.500 ;
        RECT 303.840 56.205 306.375 56.345 ;
        RECT 303.840 56.160 304.130 56.205 ;
        RECT 285.460 55.865 286.225 56.005 ;
        RECT 285.460 55.820 285.750 55.865 ;
        RECT 285.905 55.805 286.225 55.865 ;
        RECT 294.200 55.820 294.490 56.050 ;
        RECT 307.080 56.005 307.370 56.050 ;
        RECT 307.525 56.005 307.845 56.065 ;
        RECT 307.080 55.865 307.845 56.005 ;
        RECT 307.080 55.820 307.370 55.865 ;
        RECT 307.525 55.805 307.845 55.865 ;
        RECT 308.905 55.805 309.225 56.065 ;
        RECT 263.365 55.525 276.015 55.665 ;
        RECT 276.210 55.665 276.500 55.710 ;
        RECT 278.100 55.665 278.390 55.710 ;
        RECT 281.220 55.665 281.510 55.710 ;
        RECT 300.180 55.665 300.470 55.710 ;
        RECT 276.210 55.525 281.510 55.665 ;
        RECT 263.365 55.465 263.685 55.525 ;
        RECT 276.210 55.480 276.500 55.525 ;
        RECT 278.100 55.480 278.390 55.525 ;
        RECT 281.220 55.480 281.510 55.525 ;
        RECT 281.855 55.525 300.470 55.665 ;
        RECT 223.805 55.185 236.455 55.325 ;
        RECT 223.805 55.125 224.125 55.185 ;
        RECT 239.905 55.125 240.225 55.385 ;
        RECT 241.745 55.325 242.065 55.385 ;
        RECT 243.600 55.325 243.890 55.370 ;
        RECT 241.745 55.185 243.890 55.325 ;
        RECT 241.745 55.125 242.065 55.185 ;
        RECT 243.600 55.140 243.890 55.185 ;
        RECT 250.960 55.325 251.250 55.370 ;
        RECT 257.385 55.325 257.705 55.385 ;
        RECT 250.960 55.185 257.705 55.325 ;
        RECT 250.960 55.140 251.250 55.185 ;
        RECT 257.385 55.125 257.705 55.185 ;
        RECT 269.345 55.325 269.665 55.385 ;
        RECT 281.855 55.325 281.995 55.525 ;
        RECT 300.180 55.480 300.470 55.525 ;
        RECT 303.860 55.665 304.150 55.710 ;
        RECT 306.620 55.665 306.910 55.710 ;
        RECT 308.460 55.665 308.750 55.710 ;
        RECT 303.860 55.525 308.750 55.665 ;
        RECT 303.860 55.480 304.150 55.525 ;
        RECT 306.620 55.480 306.910 55.525 ;
        RECT 308.460 55.480 308.750 55.525 ;
        RECT 269.345 55.185 281.995 55.325 ;
        RECT 269.345 55.125 269.665 55.185 ;
        RECT 291.425 55.125 291.745 55.385 ;
        RECT 162.095 54.505 311.135 54.985 ;
        RECT 181.040 54.305 181.330 54.350 ;
        RECT 183.325 54.305 183.645 54.365 ;
        RECT 181.040 54.165 183.645 54.305 ;
        RECT 181.040 54.120 181.330 54.165 ;
        RECT 183.325 54.105 183.645 54.165 ;
        RECT 185.640 54.305 185.930 54.350 ;
        RECT 187.005 54.305 187.325 54.365 ;
        RECT 185.640 54.165 187.325 54.305 ;
        RECT 185.640 54.120 185.930 54.165 ;
        RECT 187.005 54.105 187.325 54.165 ;
        RECT 187.940 54.120 188.230 54.350 ;
        RECT 202.660 54.305 202.950 54.350 ;
        RECT 203.565 54.305 203.885 54.365 ;
        RECT 202.660 54.165 203.885 54.305 ;
        RECT 202.660 54.120 202.950 54.165 ;
        RECT 166.730 53.965 167.020 54.010 ;
        RECT 168.620 53.965 168.910 54.010 ;
        RECT 171.740 53.965 172.030 54.010 ;
        RECT 166.730 53.825 172.030 53.965 ;
        RECT 166.730 53.780 167.020 53.825 ;
        RECT 168.620 53.780 168.910 53.825 ;
        RECT 171.740 53.780 172.030 53.825 ;
        RECT 174.600 53.965 174.890 54.010 ;
        RECT 175.965 53.965 176.285 54.025 ;
        RECT 183.785 53.965 184.105 54.025 ;
        RECT 174.600 53.825 176.285 53.965 ;
        RECT 174.600 53.780 174.890 53.825 ;
        RECT 175.965 53.765 176.285 53.825 ;
        RECT 181.575 53.825 184.105 53.965 ;
        RECT 167.225 53.425 167.545 53.685 ;
        RECT 173.665 53.625 173.985 53.685 ;
        RECT 176.885 53.625 177.205 53.685 ;
        RECT 178.280 53.625 178.570 53.670 ;
        RECT 173.665 53.485 178.570 53.625 ;
        RECT 173.665 53.425 173.985 53.485 ;
        RECT 176.885 53.425 177.205 53.485 ;
        RECT 178.280 53.440 178.570 53.485 ;
        RECT 165.845 53.085 166.165 53.345 ;
        RECT 166.325 53.285 166.615 53.330 ;
        RECT 168.160 53.285 168.450 53.330 ;
        RECT 171.740 53.285 172.030 53.330 ;
        RECT 166.325 53.145 172.030 53.285 ;
        RECT 166.325 53.100 166.615 53.145 ;
        RECT 168.160 53.100 168.450 53.145 ;
        RECT 171.740 53.100 172.030 53.145 ;
        RECT 172.745 53.305 173.065 53.345 ;
        RECT 172.745 53.085 173.110 53.305 ;
        RECT 177.820 53.285 178.110 53.330 ;
        RECT 180.105 53.285 180.425 53.345 ;
        RECT 181.575 53.330 181.715 53.825 ;
        RECT 183.785 53.765 184.105 53.825 ;
        RECT 184.245 53.965 184.565 54.025 ;
        RECT 186.085 53.965 186.405 54.025 ;
        RECT 188.015 53.965 188.155 54.120 ;
        RECT 203.565 54.105 203.885 54.165 ;
        RECT 206.785 54.105 207.105 54.365 ;
        RECT 213.225 54.305 213.545 54.365 ;
        RECT 213.225 54.165 218.975 54.305 ;
        RECT 213.225 54.105 213.545 54.165 ;
        RECT 184.245 53.825 188.155 53.965 ;
        RECT 188.860 53.965 189.150 54.010 ;
        RECT 194.365 53.965 194.685 54.025 ;
        RECT 188.860 53.825 194.685 53.965 ;
        RECT 184.245 53.765 184.565 53.825 ;
        RECT 186.085 53.765 186.405 53.825 ;
        RECT 188.860 53.780 189.150 53.825 ;
        RECT 190.315 53.670 190.455 53.825 ;
        RECT 194.365 53.765 194.685 53.825 ;
        RECT 198.965 53.965 199.285 54.025 ;
        RECT 198.965 53.825 205.175 53.965 ;
        RECT 198.965 53.765 199.285 53.825 ;
        RECT 190.240 53.440 190.530 53.670 ;
        RECT 192.065 53.625 192.385 53.685 ;
        RECT 190.775 53.485 192.385 53.625 ;
        RECT 177.820 53.145 180.425 53.285 ;
        RECT 177.820 53.100 178.110 53.145 ;
        RECT 180.105 53.085 180.425 53.145 ;
        RECT 181.500 53.100 181.790 53.330 ;
        RECT 182.880 53.285 183.170 53.330 ;
        RECT 186.100 53.285 186.390 53.330 ;
        RECT 187.005 53.285 187.325 53.345 ;
        RECT 187.925 53.285 188.245 53.345 ;
        RECT 190.775 53.330 190.915 53.485 ;
        RECT 192.065 53.425 192.385 53.485 ;
        RECT 192.540 53.625 192.830 53.670 ;
        RECT 192.540 53.485 199.655 53.625 ;
        RECT 192.540 53.440 192.830 53.485 ;
        RECT 190.700 53.285 190.990 53.330 ;
        RECT 182.880 53.145 187.325 53.285 ;
        RECT 182.880 53.100 183.170 53.145 ;
        RECT 186.100 53.100 186.390 53.145 ;
        RECT 187.005 53.085 187.325 53.145 ;
        RECT 187.555 53.145 190.990 53.285 ;
        RECT 172.820 52.990 173.110 53.085 ;
        RECT 169.520 52.945 170.170 52.990 ;
        RECT 172.820 52.945 173.410 52.990 ;
        RECT 169.520 52.805 173.410 52.945 ;
        RECT 169.520 52.760 170.170 52.805 ;
        RECT 173.120 52.760 173.410 52.805 ;
        RECT 177.360 52.945 177.650 52.990 ;
        RECT 180.565 52.945 180.885 53.005 ;
        RECT 177.360 52.805 180.885 52.945 ;
        RECT 177.360 52.760 177.650 52.805 ;
        RECT 180.565 52.745 180.885 52.805 ;
        RECT 183.800 52.945 184.090 52.990 ;
        RECT 187.555 52.945 187.695 53.145 ;
        RECT 187.925 53.085 188.245 53.145 ;
        RECT 190.700 53.100 190.990 53.145 ;
        RECT 191.145 53.085 191.465 53.345 ;
        RECT 191.620 53.100 191.910 53.330 ;
        RECT 193.445 53.285 193.765 53.345 ;
        RECT 198.135 53.330 198.275 53.485 ;
        RECT 193.445 53.145 197.815 53.285 ;
        RECT 191.695 52.945 191.835 53.100 ;
        RECT 193.445 53.085 193.765 53.145 ;
        RECT 183.800 52.805 187.695 52.945 ;
        RECT 188.015 52.805 191.835 52.945 ;
        RECT 183.800 52.760 184.090 52.805 ;
        RECT 175.505 52.405 175.825 52.665 ;
        RECT 184.245 52.405 184.565 52.665 ;
        RECT 184.705 52.605 185.025 52.665 ;
        RECT 188.015 52.650 188.155 52.805 ;
        RECT 193.905 52.745 194.225 53.005 ;
        RECT 197.675 52.990 197.815 53.145 ;
        RECT 198.060 53.100 198.350 53.330 ;
        RECT 198.980 53.100 199.270 53.330 ;
        RECT 199.515 53.285 199.655 53.485 ;
        RECT 199.885 53.425 200.205 53.685 ;
        RECT 205.035 53.670 205.175 53.825 ;
        RECT 204.960 53.440 205.250 53.670 ;
        RECT 205.880 53.285 206.170 53.330 ;
        RECT 199.515 53.145 206.170 53.285 ;
        RECT 205.880 53.100 206.170 53.145 ;
        RECT 197.600 52.945 197.890 52.990 ;
        RECT 198.505 52.945 198.825 53.005 ;
        RECT 197.600 52.805 198.825 52.945 ;
        RECT 197.600 52.760 197.890 52.805 ;
        RECT 198.505 52.745 198.825 52.805 ;
        RECT 199.055 52.665 199.195 53.100 ;
        RECT 203.580 52.945 203.870 52.990 ;
        RECT 204.025 52.945 204.345 53.005 ;
        RECT 203.580 52.805 204.345 52.945 ;
        RECT 203.580 52.760 203.870 52.805 ;
        RECT 204.025 52.745 204.345 52.805 ;
        RECT 204.500 52.945 204.790 52.990 ;
        RECT 206.875 52.945 207.015 54.105 ;
        RECT 218.835 54.010 218.975 54.165 ;
        RECT 221.045 54.105 221.365 54.365 ;
        RECT 238.065 54.105 238.385 54.365 ;
        RECT 252.325 54.305 252.645 54.365 ;
        RECT 262.905 54.305 263.225 54.365 ;
        RECT 288.205 54.305 288.525 54.365 ;
        RECT 252.325 54.165 263.225 54.305 ;
        RECT 252.325 54.105 252.645 54.165 ;
        RECT 262.905 54.105 263.225 54.165 ;
        RECT 264.835 54.165 288.525 54.305 ;
        RECT 210.890 53.965 211.180 54.010 ;
        RECT 212.780 53.965 213.070 54.010 ;
        RECT 215.900 53.965 216.190 54.010 ;
        RECT 210.890 53.825 216.190 53.965 ;
        RECT 210.890 53.780 211.180 53.825 ;
        RECT 212.780 53.780 213.070 53.825 ;
        RECT 215.900 53.780 216.190 53.825 ;
        RECT 218.760 53.965 219.050 54.010 ;
        RECT 246.345 53.965 246.665 54.025 ;
        RECT 264.285 53.965 264.605 54.025 ;
        RECT 218.760 53.825 240.135 53.965 ;
        RECT 218.760 53.780 219.050 53.825 ;
        RECT 211.400 53.625 211.690 53.670 ;
        RECT 211.845 53.625 212.165 53.685 ;
        RECT 211.400 53.485 212.165 53.625 ;
        RECT 211.400 53.440 211.690 53.485 ;
        RECT 211.845 53.425 212.165 53.485 ;
        RECT 225.660 53.625 225.950 53.670 ;
        RECT 227.485 53.625 227.805 53.685 ;
        RECT 239.995 53.670 240.135 53.825 ;
        RECT 246.345 53.825 264.605 53.965 ;
        RECT 246.345 53.765 246.665 53.825 ;
        RECT 264.285 53.765 264.605 53.825 ;
        RECT 225.660 53.485 227.805 53.625 ;
        RECT 225.660 53.440 225.950 53.485 ;
        RECT 227.485 53.425 227.805 53.485 ;
        RECT 239.920 53.440 240.210 53.670 ;
        RECT 240.380 53.625 240.670 53.670 ;
        RECT 242.220 53.625 242.510 53.670 ;
        RECT 240.380 53.485 242.510 53.625 ;
        RECT 240.380 53.440 240.670 53.485 ;
        RECT 242.220 53.440 242.510 53.485 ;
        RECT 252.785 53.625 253.105 53.685 ;
        RECT 263.840 53.625 264.130 53.670 ;
        RECT 252.785 53.485 264.130 53.625 ;
        RECT 252.785 53.425 253.105 53.485 ;
        RECT 263.840 53.440 264.130 53.485 ;
        RECT 210.020 53.100 210.310 53.330 ;
        RECT 210.485 53.285 210.775 53.330 ;
        RECT 212.320 53.285 212.610 53.330 ;
        RECT 215.900 53.285 216.190 53.330 ;
        RECT 210.485 53.145 216.190 53.285 ;
        RECT 210.485 53.100 210.775 53.145 ;
        RECT 212.320 53.100 212.610 53.145 ;
        RECT 215.900 53.100 216.190 53.145 ;
        RECT 210.095 52.945 210.235 53.100 ;
        RECT 216.980 52.990 217.270 53.305 ;
        RECT 218.745 53.085 219.065 53.345 ;
        RECT 219.205 53.285 219.525 53.345 ;
        RECT 219.205 53.145 220.815 53.285 ;
        RECT 219.205 53.085 219.525 53.145 ;
        RECT 204.500 52.805 207.015 52.945 ;
        RECT 207.335 52.805 210.235 52.945 ;
        RECT 213.680 52.945 214.330 52.990 ;
        RECT 216.980 52.945 217.570 52.990 ;
        RECT 218.835 52.945 218.975 53.085 ;
        RECT 220.140 52.945 220.430 52.990 ;
        RECT 213.680 52.805 218.515 52.945 ;
        RECT 218.835 52.805 220.430 52.945 ;
        RECT 220.675 52.945 220.815 53.145 ;
        RECT 221.505 53.085 221.825 53.345 ;
        RECT 227.945 53.085 228.265 53.345 ;
        RECT 239.000 53.285 239.290 53.330 ;
        RECT 239.000 53.145 240.595 53.285 ;
        RECT 239.000 53.100 239.290 53.145 ;
        RECT 225.645 52.945 225.965 53.005 ;
        RECT 220.675 52.805 225.965 52.945 ;
        RECT 204.500 52.760 204.790 52.805 ;
        RECT 187.940 52.605 188.230 52.650 ;
        RECT 184.705 52.465 188.230 52.605 ;
        RECT 184.705 52.405 185.025 52.465 ;
        RECT 187.940 52.420 188.230 52.465 ;
        RECT 194.825 52.605 195.145 52.665 ;
        RECT 198.965 52.605 199.285 52.665 ;
        RECT 194.825 52.465 199.285 52.605 ;
        RECT 194.825 52.405 195.145 52.465 ;
        RECT 198.965 52.405 199.285 52.465 ;
        RECT 200.805 52.605 201.125 52.665 ;
        RECT 207.335 52.605 207.475 52.805 ;
        RECT 213.680 52.760 214.330 52.805 ;
        RECT 217.280 52.760 217.570 52.805 ;
        RECT 200.805 52.465 207.475 52.605 ;
        RECT 211.385 52.605 211.705 52.665 ;
        RECT 218.375 52.605 218.515 52.805 ;
        RECT 220.140 52.760 220.430 52.805 ;
        RECT 225.645 52.745 225.965 52.805 ;
        RECT 222.885 52.605 223.205 52.665 ;
        RECT 211.385 52.465 223.205 52.605 ;
        RECT 240.455 52.605 240.595 53.145 ;
        RECT 240.840 53.100 241.130 53.330 ;
        RECT 240.915 52.945 241.055 53.100 ;
        RECT 241.745 53.085 242.065 53.345 ;
        RECT 244.965 53.085 245.285 53.345 ;
        RECT 245.900 53.100 246.190 53.330 ;
        RECT 258.305 53.285 258.625 53.345 ;
        RECT 263.380 53.285 263.670 53.330 ;
        RECT 264.835 53.285 264.975 54.165 ;
        RECT 288.205 54.105 288.525 54.165 ;
        RECT 297.865 54.305 298.185 54.365 ;
        RECT 302.020 54.305 302.310 54.350 ;
        RECT 297.865 54.165 302.310 54.305 ;
        RECT 297.865 54.105 298.185 54.165 ;
        RECT 302.020 54.120 302.310 54.165 ;
        RECT 307.525 54.105 307.845 54.365 ;
        RECT 280.385 53.965 280.705 54.025 ;
        RECT 269.665 53.825 280.705 53.965 ;
        RECT 269.665 53.625 269.805 53.825 ;
        RECT 280.385 53.765 280.705 53.825 ;
        RECT 281.420 53.965 281.710 54.010 ;
        RECT 284.540 53.965 284.830 54.010 ;
        RECT 286.430 53.965 286.720 54.010 ;
        RECT 281.420 53.825 286.720 53.965 ;
        RECT 281.420 53.780 281.710 53.825 ;
        RECT 284.540 53.780 284.830 53.825 ;
        RECT 286.430 53.780 286.720 53.825 ;
        RECT 291.885 53.965 292.205 54.025 ;
        RECT 308.460 53.965 308.750 54.010 ;
        RECT 291.885 53.825 308.750 53.965 ;
        RECT 291.885 53.765 292.205 53.825 ;
        RECT 308.460 53.780 308.750 53.825 ;
        RECT 268.975 53.485 269.805 53.625 ;
        RECT 275.325 53.625 275.645 53.685 ;
        RECT 285.905 53.625 286.225 53.685 ;
        RECT 275.325 53.485 286.225 53.625 ;
        RECT 258.305 53.145 264.975 53.285 ;
        RECT 242.665 52.945 242.985 53.005 ;
        RECT 240.915 52.805 242.985 52.945 ;
        RECT 242.665 52.745 242.985 52.805 ;
        RECT 244.505 52.945 244.825 53.005 ;
        RECT 245.975 52.945 246.115 53.100 ;
        RECT 258.305 53.085 258.625 53.145 ;
        RECT 263.380 53.100 263.670 53.145 ;
        RECT 266.585 53.085 266.905 53.345 ;
        RECT 267.505 53.085 267.825 53.345 ;
        RECT 267.965 53.285 268.285 53.345 ;
        RECT 268.975 53.330 269.115 53.485 ;
        RECT 275.325 53.425 275.645 53.485 ;
        RECT 267.965 53.145 268.480 53.285 ;
        RECT 267.965 53.085 268.285 53.145 ;
        RECT 268.900 53.100 269.190 53.330 ;
        RECT 269.345 53.085 269.665 53.345 ;
        RECT 276.335 53.330 276.475 53.485 ;
        RECT 285.905 53.425 286.225 53.485 ;
        RECT 287.300 53.625 287.590 53.670 ;
        RECT 290.505 53.625 290.825 53.685 ;
        RECT 291.440 53.625 291.730 53.670 ;
        RECT 287.300 53.485 291.730 53.625 ;
        RECT 287.300 53.440 287.590 53.485 ;
        RECT 290.505 53.425 290.825 53.485 ;
        RECT 291.440 53.440 291.730 53.485 ;
        RECT 269.845 53.100 270.135 53.330 ;
        RECT 276.260 53.100 276.550 53.330 ;
        RECT 244.505 52.805 246.115 52.945 ;
        RECT 254.165 52.945 254.485 53.005 ;
        RECT 254.640 52.945 254.930 52.990 ;
        RECT 255.545 52.945 255.865 53.005 ;
        RECT 254.165 52.805 255.865 52.945 ;
        RECT 244.505 52.745 244.825 52.805 ;
        RECT 254.165 52.745 254.485 52.805 ;
        RECT 254.640 52.760 254.930 52.805 ;
        RECT 255.545 52.745 255.865 52.805 ;
        RECT 258.765 52.945 259.085 53.005 ;
        RECT 259.240 52.945 259.530 52.990 ;
        RECT 258.765 52.805 259.530 52.945 ;
        RECT 258.765 52.745 259.085 52.805 ;
        RECT 259.240 52.760 259.530 52.805 ;
        RECT 262.905 52.945 263.225 53.005 ;
        RECT 269.435 52.945 269.575 53.085 ;
        RECT 262.905 52.805 269.575 52.945 ;
        RECT 262.905 52.745 263.225 52.805 ;
        RECT 241.285 52.605 241.605 52.665 ;
        RECT 240.455 52.465 241.605 52.605 ;
        RECT 200.805 52.405 201.125 52.465 ;
        RECT 211.385 52.405 211.705 52.465 ;
        RECT 222.885 52.405 223.205 52.465 ;
        RECT 241.285 52.405 241.605 52.465 ;
        RECT 249.105 52.405 249.425 52.665 ;
        RECT 257.845 52.605 258.165 52.665 ;
        RECT 269.920 52.605 270.060 53.100 ;
        RECT 278.085 52.945 278.405 53.005 ;
        RECT 280.340 52.990 280.630 53.305 ;
        RECT 281.420 53.285 281.710 53.330 ;
        RECT 285.000 53.285 285.290 53.330 ;
        RECT 286.835 53.285 287.125 53.330 ;
        RECT 281.420 53.145 287.125 53.285 ;
        RECT 281.420 53.100 281.710 53.145 ;
        RECT 285.000 53.100 285.290 53.145 ;
        RECT 286.835 53.100 287.125 53.145 ;
        RECT 287.760 53.285 288.050 53.330 ;
        RECT 288.205 53.285 288.525 53.345 ;
        RECT 287.760 53.145 288.525 53.285 ;
        RECT 287.760 53.100 288.050 53.145 ;
        RECT 288.205 53.085 288.525 53.145 ;
        RECT 300.165 53.285 300.485 53.345 ;
        RECT 304.320 53.285 304.610 53.330 ;
        RECT 300.165 53.145 304.610 53.285 ;
        RECT 300.165 53.085 300.485 53.145 ;
        RECT 304.320 53.100 304.610 53.145 ;
        RECT 309.365 53.085 309.685 53.345 ;
        RECT 280.040 52.945 280.630 52.990 ;
        RECT 283.280 52.945 283.930 52.990 ;
        RECT 278.085 52.805 283.930 52.945 ;
        RECT 278.085 52.745 278.405 52.805 ;
        RECT 280.040 52.760 280.330 52.805 ;
        RECT 283.280 52.760 283.930 52.805 ;
        RECT 285.920 52.945 286.210 52.990 ;
        RECT 291.425 52.945 291.745 53.005 ;
        RECT 285.920 52.805 291.745 52.945 ;
        RECT 285.920 52.760 286.210 52.805 ;
        RECT 291.425 52.745 291.745 52.805 ;
        RECT 294.185 52.945 294.505 53.005 ;
        RECT 301.560 52.945 301.850 52.990 ;
        RECT 303.845 52.945 304.165 53.005 ;
        RECT 294.185 52.805 304.165 52.945 ;
        RECT 294.185 52.745 294.505 52.805 ;
        RECT 301.560 52.760 301.850 52.805 ;
        RECT 303.845 52.745 304.165 52.805 ;
        RECT 257.845 52.465 270.060 52.605 ;
        RECT 257.845 52.405 258.165 52.465 ;
        RECT 270.725 52.405 271.045 52.665 ;
        RECT 278.545 52.405 278.865 52.665 ;
        RECT 162.095 51.785 311.135 52.265 ;
        RECT 175.505 51.585 175.825 51.645 ;
        RECT 167.315 51.445 175.825 51.585 ;
        RECT 167.315 51.290 167.455 51.445 ;
        RECT 175.505 51.385 175.825 51.445 ;
        RECT 176.885 51.585 177.205 51.645 ;
        RECT 184.260 51.585 184.550 51.630 ;
        RECT 176.885 51.445 184.550 51.585 ;
        RECT 176.885 51.385 177.205 51.445 ;
        RECT 184.260 51.400 184.550 51.445 ;
        RECT 186.100 51.585 186.390 51.630 ;
        RECT 187.465 51.585 187.785 51.645 ;
        RECT 194.825 51.585 195.145 51.645 ;
        RECT 200.805 51.585 201.125 51.645 ;
        RECT 214.145 51.585 214.465 51.645 ;
        RECT 221.965 51.585 222.285 51.645 ;
        RECT 225.185 51.585 225.505 51.645 ;
        RECT 260.605 51.585 260.925 51.645 ;
        RECT 264.760 51.585 265.050 51.630 ;
        RECT 266.585 51.585 266.905 51.645 ;
        RECT 276.705 51.585 277.025 51.645 ;
        RECT 300.165 51.630 300.485 51.645 ;
        RECT 186.100 51.445 195.145 51.585 ;
        RECT 186.100 51.400 186.390 51.445 ;
        RECT 187.465 51.385 187.785 51.445 ;
        RECT 194.825 51.385 195.145 51.445 ;
        RECT 195.375 51.445 201.125 51.585 ;
        RECT 178.725 51.290 179.045 51.305 ;
        RECT 167.240 51.060 167.530 51.290 ;
        RECT 169.520 51.245 170.170 51.290 ;
        RECT 173.120 51.245 173.410 51.290 ;
        RECT 178.720 51.245 179.370 51.290 ;
        RECT 182.320 51.245 182.610 51.290 ;
        RECT 169.520 51.105 182.610 51.245 ;
        RECT 169.520 51.060 170.170 51.105 ;
        RECT 172.820 51.060 173.410 51.105 ;
        RECT 178.720 51.060 179.370 51.105 ;
        RECT 182.020 51.060 182.610 51.105 ;
        RECT 184.705 51.245 185.025 51.305 ;
        RECT 191.160 51.245 191.450 51.290 ;
        RECT 184.705 51.105 191.450 51.245 ;
        RECT 172.820 50.965 173.205 51.060 ;
        RECT 178.725 51.045 179.045 51.060 ;
        RECT 166.325 50.905 166.615 50.950 ;
        RECT 168.160 50.905 168.450 50.950 ;
        RECT 171.740 50.905 172.030 50.950 ;
        RECT 166.325 50.765 172.030 50.905 ;
        RECT 166.325 50.720 166.615 50.765 ;
        RECT 168.160 50.720 168.450 50.765 ;
        RECT 171.740 50.720 172.030 50.765 ;
        RECT 172.745 50.765 173.205 50.965 ;
        RECT 172.745 50.745 173.110 50.765 ;
        RECT 172.745 50.705 173.065 50.745 ;
        RECT 175.045 50.705 175.365 50.965 ;
        RECT 175.525 50.905 175.815 50.950 ;
        RECT 177.360 50.905 177.650 50.950 ;
        RECT 180.940 50.905 181.230 50.950 ;
        RECT 175.525 50.765 181.230 50.905 ;
        RECT 175.525 50.720 175.815 50.765 ;
        RECT 177.360 50.720 177.650 50.765 ;
        RECT 180.940 50.720 181.230 50.765 ;
        RECT 182.020 50.745 182.310 51.060 ;
        RECT 184.705 51.045 185.025 51.105 ;
        RECT 191.160 51.060 191.450 51.105 ;
        RECT 192.080 51.245 192.370 51.290 ;
        RECT 192.985 51.245 193.305 51.305 ;
        RECT 192.080 51.105 193.305 51.245 ;
        RECT 192.080 51.060 192.370 51.105 ;
        RECT 192.985 51.045 193.305 51.105 ;
        RECT 190.240 50.720 190.530 50.950 ;
        RECT 165.845 50.365 166.165 50.625 ;
        RECT 174.585 50.365 174.905 50.625 ;
        RECT 176.425 50.365 176.745 50.625 ;
        RECT 183.785 50.365 184.105 50.625 ;
        RECT 185.055 50.380 185.345 50.610 ;
        RECT 166.730 50.225 167.020 50.270 ;
        RECT 168.620 50.225 168.910 50.270 ;
        RECT 171.740 50.225 172.030 50.270 ;
        RECT 166.730 50.085 172.030 50.225 ;
        RECT 166.730 50.040 167.020 50.085 ;
        RECT 168.620 50.040 168.910 50.085 ;
        RECT 171.740 50.040 172.030 50.085 ;
        RECT 175.930 50.225 176.220 50.270 ;
        RECT 177.820 50.225 178.110 50.270 ;
        RECT 180.940 50.225 181.230 50.270 ;
        RECT 175.930 50.085 181.230 50.225 ;
        RECT 185.130 50.225 185.270 50.380 ;
        RECT 185.625 50.365 185.945 50.625 ;
        RECT 187.480 50.565 187.770 50.610 ;
        RECT 187.925 50.565 188.245 50.625 ;
        RECT 190.315 50.565 190.455 50.720 ;
        RECT 190.685 50.705 191.005 50.965 ;
        RECT 194.380 50.905 194.670 50.950 ;
        RECT 195.375 50.905 195.515 51.445 ;
        RECT 200.805 51.385 201.125 51.445 ;
        RECT 204.575 51.445 214.465 51.585 ;
        RECT 198.045 51.245 198.365 51.305 ;
        RECT 198.960 51.245 199.610 51.290 ;
        RECT 202.560 51.245 202.850 51.290 ;
        RECT 198.045 51.105 202.850 51.245 ;
        RECT 198.045 51.045 198.365 51.105 ;
        RECT 198.960 51.060 199.610 51.105 ;
        RECT 202.260 51.060 202.850 51.105 ;
        RECT 194.380 50.765 195.515 50.905 ;
        RECT 195.765 50.905 196.055 50.950 ;
        RECT 197.600 50.905 197.890 50.950 ;
        RECT 201.180 50.905 201.470 50.950 ;
        RECT 195.765 50.765 201.470 50.905 ;
        RECT 194.380 50.720 194.670 50.765 ;
        RECT 195.765 50.720 196.055 50.765 ;
        RECT 197.600 50.720 197.890 50.765 ;
        RECT 201.180 50.720 201.470 50.765 ;
        RECT 202.260 50.745 202.550 51.060 ;
        RECT 204.575 50.950 204.715 51.445 ;
        RECT 214.145 51.385 214.465 51.445 ;
        RECT 214.695 51.445 223.575 51.585 ;
        RECT 205.880 51.245 206.170 51.290 ;
        RECT 207.245 51.245 207.565 51.305 ;
        RECT 205.880 51.105 207.565 51.245 ;
        RECT 205.880 51.060 206.170 51.105 ;
        RECT 207.245 51.045 207.565 51.105 ;
        RECT 208.160 51.245 208.810 51.290 ;
        RECT 211.760 51.245 212.050 51.290 ;
        RECT 214.695 51.245 214.835 51.445 ;
        RECT 221.965 51.385 222.285 51.445 ;
        RECT 208.160 51.105 212.050 51.245 ;
        RECT 208.160 51.060 208.810 51.105 ;
        RECT 211.460 51.060 212.050 51.105 ;
        RECT 212.395 51.105 214.835 51.245 ;
        RECT 215.065 51.245 215.385 51.305 ;
        RECT 223.435 51.290 223.575 51.445 ;
        RECT 225.185 51.445 248.415 51.585 ;
        RECT 225.185 51.385 225.505 51.445 ;
        RECT 215.540 51.245 215.830 51.290 ;
        RECT 215.065 51.105 215.830 51.245 ;
        RECT 211.460 50.965 211.750 51.060 ;
        RECT 204.500 50.720 204.790 50.950 ;
        RECT 204.965 50.905 205.255 50.950 ;
        RECT 206.800 50.905 207.090 50.950 ;
        RECT 210.380 50.905 210.670 50.950 ;
        RECT 204.965 50.765 210.670 50.905 ;
        RECT 204.965 50.720 205.255 50.765 ;
        RECT 206.800 50.720 207.090 50.765 ;
        RECT 210.380 50.720 210.670 50.765 ;
        RECT 211.385 50.745 211.750 50.965 ;
        RECT 211.385 50.705 211.705 50.745 ;
        RECT 187.480 50.425 190.455 50.565 ;
        RECT 193.905 50.565 194.225 50.625 ;
        RECT 195.300 50.565 195.590 50.610 ;
        RECT 193.905 50.425 195.590 50.565 ;
        RECT 187.480 50.380 187.770 50.425 ;
        RECT 187.925 50.365 188.245 50.425 ;
        RECT 193.905 50.365 194.225 50.425 ;
        RECT 195.300 50.380 195.590 50.425 ;
        RECT 198.505 50.565 198.825 50.625 ;
        RECT 198.505 50.425 204.715 50.565 ;
        RECT 198.505 50.365 198.825 50.425 ;
        RECT 187.005 50.225 187.325 50.285 ;
        RECT 189.320 50.225 189.610 50.270 ;
        RECT 190.225 50.225 190.545 50.285 ;
        RECT 185.130 50.085 190.545 50.225 ;
        RECT 175.930 50.040 176.220 50.085 ;
        RECT 177.820 50.040 178.110 50.085 ;
        RECT 180.940 50.040 181.230 50.085 ;
        RECT 187.005 50.025 187.325 50.085 ;
        RECT 189.320 50.040 189.610 50.085 ;
        RECT 190.225 50.025 190.545 50.085 ;
        RECT 196.170 50.225 196.460 50.270 ;
        RECT 198.060 50.225 198.350 50.270 ;
        RECT 201.180 50.225 201.470 50.270 ;
        RECT 196.170 50.085 201.470 50.225 ;
        RECT 196.170 50.040 196.460 50.085 ;
        RECT 198.060 50.040 198.350 50.085 ;
        RECT 201.180 50.040 201.470 50.085 ;
        RECT 204.025 50.025 204.345 50.285 ;
        RECT 196.615 49.885 196.905 49.930 ;
        RECT 201.725 49.885 202.045 49.945 ;
        RECT 196.615 49.745 202.045 49.885 ;
        RECT 204.575 49.885 204.715 50.425 ;
        RECT 205.370 50.225 205.660 50.270 ;
        RECT 207.260 50.225 207.550 50.270 ;
        RECT 210.380 50.225 210.670 50.270 ;
        RECT 205.370 50.085 210.670 50.225 ;
        RECT 205.370 50.040 205.660 50.085 ;
        RECT 207.260 50.040 207.550 50.085 ;
        RECT 210.380 50.040 210.670 50.085 ;
        RECT 212.395 49.885 212.535 51.105 ;
        RECT 215.065 51.045 215.385 51.105 ;
        RECT 215.540 51.060 215.830 51.105 ;
        RECT 217.820 51.245 218.470 51.290 ;
        RECT 221.420 51.245 221.710 51.290 ;
        RECT 217.820 51.105 221.710 51.245 ;
        RECT 217.820 51.060 218.470 51.105 ;
        RECT 221.120 51.060 221.710 51.105 ;
        RECT 223.360 51.060 223.650 51.290 ;
        RECT 233.920 51.245 234.570 51.290 ;
        RECT 237.520 51.245 237.810 51.290 ;
        RECT 233.920 51.105 237.810 51.245 ;
        RECT 233.920 51.060 234.570 51.105 ;
        RECT 237.220 51.060 237.810 51.105 ;
        RECT 239.445 51.245 239.765 51.305 ;
        RECT 246.345 51.245 246.665 51.305 ;
        RECT 239.445 51.105 241.975 51.245 ;
        RECT 214.625 50.905 214.915 50.950 ;
        RECT 216.460 50.905 216.750 50.950 ;
        RECT 220.040 50.905 220.330 50.950 ;
        RECT 214.625 50.765 220.330 50.905 ;
        RECT 214.625 50.720 214.915 50.765 ;
        RECT 216.460 50.720 216.750 50.765 ;
        RECT 220.040 50.720 220.330 50.765 ;
        RECT 221.120 50.905 221.410 51.060 ;
        RECT 237.220 50.965 237.510 51.060 ;
        RECT 239.445 51.045 239.765 51.105 ;
        RECT 222.885 50.905 223.205 50.965 ;
        RECT 226.105 50.905 226.425 50.965 ;
        RECT 221.120 50.765 226.425 50.905 ;
        RECT 221.120 50.745 221.410 50.765 ;
        RECT 222.885 50.705 223.205 50.765 ;
        RECT 226.105 50.705 226.425 50.765 ;
        RECT 230.725 50.905 231.015 50.950 ;
        RECT 232.560 50.905 232.850 50.950 ;
        RECT 236.140 50.905 236.430 50.950 ;
        RECT 230.725 50.765 236.430 50.905 ;
        RECT 230.725 50.720 231.015 50.765 ;
        RECT 232.560 50.720 232.850 50.765 ;
        RECT 236.140 50.720 236.430 50.765 ;
        RECT 237.145 50.745 237.510 50.965 ;
        RECT 240.840 50.905 241.130 50.950 ;
        RECT 241.285 50.905 241.605 50.965 ;
        RECT 241.835 50.950 241.975 51.105 ;
        RECT 242.755 51.105 246.665 51.245 ;
        RECT 242.755 50.965 242.895 51.105 ;
        RECT 246.345 51.045 246.665 51.105 ;
        RECT 240.840 50.765 241.605 50.905 ;
        RECT 237.145 50.705 237.465 50.745 ;
        RECT 240.840 50.720 241.130 50.765 ;
        RECT 241.285 50.705 241.605 50.765 ;
        RECT 241.760 50.720 242.050 50.950 ;
        RECT 242.665 50.705 242.985 50.965 ;
        RECT 243.125 50.905 243.445 50.965 ;
        RECT 243.600 50.905 243.890 50.950 ;
        RECT 247.265 50.905 247.585 50.965 ;
        RECT 243.125 50.765 243.890 50.905 ;
        RECT 243.125 50.705 243.445 50.765 ;
        RECT 243.600 50.720 243.890 50.765 ;
        RECT 244.720 50.765 247.585 50.905 ;
        RECT 213.240 50.565 213.530 50.610 ;
        RECT 213.685 50.565 214.005 50.625 ;
        RECT 213.240 50.425 214.005 50.565 ;
        RECT 213.240 50.380 213.530 50.425 ;
        RECT 213.685 50.365 214.005 50.425 ;
        RECT 214.145 50.365 214.465 50.625 ;
        RECT 227.500 50.565 227.790 50.610 ;
        RECT 227.945 50.565 228.265 50.625 ;
        RECT 230.260 50.565 230.550 50.610 ;
        RECT 227.500 50.425 230.550 50.565 ;
        RECT 227.500 50.380 227.790 50.425 ;
        RECT 227.945 50.365 228.265 50.425 ;
        RECT 230.260 50.380 230.550 50.425 ;
        RECT 231.625 50.365 231.945 50.625 ;
        RECT 232.085 50.565 232.405 50.625 ;
        RECT 239.920 50.565 240.210 50.610 ;
        RECT 232.085 50.425 240.210 50.565 ;
        RECT 232.085 50.365 232.405 50.425 ;
        RECT 239.920 50.380 240.210 50.425 ;
        RECT 242.220 50.565 242.510 50.610 ;
        RECT 244.720 50.565 244.860 50.765 ;
        RECT 247.265 50.705 247.585 50.765 ;
        RECT 247.725 50.705 248.045 50.965 ;
        RECT 248.275 50.905 248.415 51.445 ;
        RECT 260.605 51.445 264.055 51.585 ;
        RECT 260.605 51.385 260.925 51.445 ;
        RECT 256.005 51.245 256.325 51.305 ;
        RECT 250.575 51.105 256.325 51.245 ;
        RECT 248.660 50.905 248.950 50.950 ;
        RECT 248.275 50.765 248.950 50.905 ;
        RECT 248.660 50.720 248.950 50.765 ;
        RECT 249.105 50.705 249.425 50.965 ;
        RECT 250.575 50.950 250.715 51.105 ;
        RECT 256.005 51.045 256.325 51.105 ;
        RECT 257.385 51.045 257.705 51.305 ;
        RECT 259.680 51.245 260.330 51.290 ;
        RECT 263.280 51.245 263.570 51.290 ;
        RECT 263.915 51.245 264.055 51.445 ;
        RECT 264.760 51.445 266.905 51.585 ;
        RECT 264.760 51.400 265.050 51.445 ;
        RECT 266.585 51.385 266.905 51.445 ;
        RECT 268.975 51.445 277.025 51.585 ;
        RECT 268.975 51.245 269.115 51.445 ;
        RECT 276.705 51.385 277.025 51.445 ;
        RECT 299.950 51.400 300.485 51.630 ;
        RECT 300.165 51.385 300.485 51.400 ;
        RECT 259.680 51.105 269.115 51.245 ;
        RECT 269.360 51.245 269.650 51.290 ;
        RECT 270.725 51.245 271.045 51.305 ;
        RECT 269.360 51.105 271.045 51.245 ;
        RECT 259.680 51.060 260.330 51.105 ;
        RECT 262.980 51.060 263.570 51.105 ;
        RECT 269.360 51.060 269.650 51.105 ;
        RECT 249.580 50.720 249.870 50.950 ;
        RECT 250.500 50.720 250.790 50.950 ;
        RECT 256.485 50.905 256.775 50.950 ;
        RECT 258.320 50.905 258.610 50.950 ;
        RECT 261.900 50.905 262.190 50.950 ;
        RECT 251.035 50.765 254.395 50.905 ;
        RECT 242.220 50.425 244.860 50.565 ;
        RECT 246.345 50.565 246.665 50.625 ;
        RECT 249.655 50.565 249.795 50.720 ;
        RECT 251.035 50.565 251.175 50.765 ;
        RECT 246.345 50.425 251.175 50.565 ;
        RECT 242.220 50.380 242.510 50.425 ;
        RECT 246.345 50.365 246.665 50.425 ;
        RECT 253.720 50.380 254.010 50.610 ;
        RECT 215.030 50.225 215.320 50.270 ;
        RECT 216.920 50.225 217.210 50.270 ;
        RECT 220.040 50.225 220.330 50.270 ;
        RECT 231.130 50.225 231.420 50.270 ;
        RECT 233.020 50.225 233.310 50.270 ;
        RECT 236.140 50.225 236.430 50.270 ;
        RECT 215.030 50.085 220.330 50.225 ;
        RECT 215.030 50.040 215.320 50.085 ;
        RECT 216.920 50.040 217.210 50.085 ;
        RECT 220.040 50.040 220.330 50.085 ;
        RECT 221.365 50.085 230.935 50.225 ;
        RECT 204.575 49.745 212.535 49.885 ;
        RECT 215.525 49.885 215.845 49.945 ;
        RECT 221.365 49.885 221.505 50.085 ;
        RECT 215.525 49.745 221.505 49.885 ;
        RECT 196.615 49.700 196.905 49.745 ;
        RECT 201.725 49.685 202.045 49.745 ;
        RECT 215.525 49.685 215.845 49.745 ;
        RECT 222.885 49.685 223.205 49.945 ;
        RECT 230.795 49.885 230.935 50.085 ;
        RECT 231.130 50.085 236.430 50.225 ;
        RECT 231.130 50.040 231.420 50.085 ;
        RECT 233.020 50.040 233.310 50.085 ;
        RECT 236.140 50.040 236.430 50.085 ;
        RECT 246.820 50.225 247.110 50.270 ;
        RECT 253.795 50.225 253.935 50.380 ;
        RECT 246.820 50.085 253.935 50.225 ;
        RECT 246.820 50.040 247.110 50.085 ;
        RECT 239.000 49.885 239.290 49.930 ;
        RECT 244.965 49.885 245.285 49.945 ;
        RECT 230.795 49.745 245.285 49.885 ;
        RECT 239.000 49.700 239.290 49.745 ;
        RECT 244.965 49.685 245.285 49.745 ;
        RECT 249.565 49.885 249.885 49.945 ;
        RECT 250.960 49.885 251.250 49.930 ;
        RECT 249.565 49.745 251.250 49.885 ;
        RECT 254.255 49.885 254.395 50.765 ;
        RECT 256.485 50.765 262.190 50.905 ;
        RECT 256.485 50.720 256.775 50.765 ;
        RECT 258.320 50.720 258.610 50.765 ;
        RECT 261.900 50.720 262.190 50.765 ;
        RECT 262.980 50.745 263.270 51.060 ;
        RECT 270.725 51.045 271.045 51.105 ;
        RECT 271.640 51.245 272.290 51.290 ;
        RECT 275.240 51.245 275.530 51.290 ;
        RECT 278.085 51.245 278.405 51.305 ;
        RECT 278.660 51.245 278.950 51.290 ;
        RECT 281.900 51.245 282.550 51.290 ;
        RECT 271.640 51.105 282.550 51.245 ;
        RECT 271.640 51.060 272.290 51.105 ;
        RECT 274.940 51.060 275.530 51.105 ;
        RECT 268.445 50.905 268.735 50.950 ;
        RECT 270.280 50.905 270.570 50.950 ;
        RECT 273.860 50.905 274.150 50.950 ;
        RECT 268.445 50.765 274.150 50.905 ;
        RECT 268.445 50.720 268.735 50.765 ;
        RECT 270.280 50.720 270.570 50.765 ;
        RECT 273.860 50.720 274.150 50.765 ;
        RECT 274.940 50.745 275.230 51.060 ;
        RECT 278.085 51.045 278.405 51.105 ;
        RECT 278.660 51.060 279.250 51.105 ;
        RECT 281.900 51.060 282.550 51.105 ;
        RECT 284.540 51.245 284.830 51.290 ;
        RECT 286.380 51.245 286.670 51.290 ;
        RECT 284.540 51.105 286.670 51.245 ;
        RECT 284.540 51.060 284.830 51.105 ;
        RECT 286.380 51.060 286.670 51.105 ;
        RECT 297.865 51.245 298.185 51.305 ;
        RECT 301.955 51.245 302.245 51.290 ;
        RECT 305.215 51.245 305.505 51.290 ;
        RECT 297.865 51.105 305.505 51.245 ;
        RECT 278.960 50.745 279.250 51.060 ;
        RECT 297.865 51.045 298.185 51.105 ;
        RECT 301.955 51.060 302.245 51.105 ;
        RECT 305.215 51.060 305.505 51.105 ;
        RECT 306.135 51.245 306.425 51.290 ;
        RECT 307.995 51.245 308.285 51.290 ;
        RECT 306.135 51.105 308.285 51.245 ;
        RECT 306.135 51.060 306.425 51.105 ;
        RECT 307.995 51.060 308.285 51.105 ;
        RECT 280.040 50.905 280.330 50.950 ;
        RECT 283.620 50.905 283.910 50.950 ;
        RECT 285.455 50.905 285.745 50.950 ;
        RECT 280.040 50.765 285.745 50.905 ;
        RECT 280.040 50.720 280.330 50.765 ;
        RECT 283.620 50.720 283.910 50.765 ;
        RECT 285.455 50.720 285.745 50.765 ;
        RECT 290.505 50.905 290.825 50.965 ;
        RECT 291.900 50.905 292.190 50.950 ;
        RECT 290.505 50.765 292.190 50.905 ;
        RECT 290.505 50.705 290.825 50.765 ;
        RECT 291.900 50.720 292.190 50.765 ;
        RECT 303.815 50.905 304.105 50.950 ;
        RECT 306.135 50.905 306.350 51.060 ;
        RECT 303.815 50.765 306.350 50.905 ;
        RECT 307.080 50.905 307.370 50.950 ;
        RECT 308.445 50.905 308.765 50.965 ;
        RECT 307.080 50.765 308.765 50.905 ;
        RECT 303.815 50.720 304.105 50.765 ;
        RECT 307.080 50.720 307.370 50.765 ;
        RECT 308.445 50.705 308.765 50.765 ;
        RECT 308.905 50.705 309.225 50.965 ;
        RECT 255.545 50.565 255.865 50.625 ;
        RECT 256.020 50.565 256.310 50.610 ;
        RECT 255.545 50.425 256.310 50.565 ;
        RECT 255.545 50.365 255.865 50.425 ;
        RECT 256.020 50.380 256.310 50.425 ;
        RECT 267.980 50.380 268.270 50.610 ;
        RECT 256.890 50.225 257.180 50.270 ;
        RECT 258.780 50.225 259.070 50.270 ;
        RECT 261.900 50.225 262.190 50.270 ;
        RECT 256.890 50.085 262.190 50.225 ;
        RECT 256.890 50.040 257.180 50.085 ;
        RECT 258.780 50.040 259.070 50.085 ;
        RECT 261.900 50.040 262.190 50.085 ;
        RECT 260.145 49.885 260.465 49.945 ;
        RECT 254.255 49.745 260.465 49.885 ;
        RECT 268.055 49.885 268.195 50.380 ;
        RECT 285.905 50.365 286.225 50.625 ;
        RECT 286.825 50.565 287.145 50.625 ;
        RECT 289.140 50.565 289.430 50.610 ;
        RECT 286.825 50.425 289.430 50.565 ;
        RECT 286.825 50.365 287.145 50.425 ;
        RECT 289.140 50.380 289.430 50.425 ;
        RECT 268.850 50.225 269.140 50.270 ;
        RECT 270.740 50.225 271.030 50.270 ;
        RECT 273.860 50.225 274.150 50.270 ;
        RECT 268.850 50.085 274.150 50.225 ;
        RECT 268.850 50.040 269.140 50.085 ;
        RECT 270.740 50.040 271.030 50.085 ;
        RECT 273.860 50.040 274.150 50.085 ;
        RECT 276.720 50.225 277.010 50.270 ;
        RECT 279.005 50.225 279.325 50.285 ;
        RECT 276.720 50.085 279.325 50.225 ;
        RECT 276.720 50.040 277.010 50.085 ;
        RECT 279.005 50.025 279.325 50.085 ;
        RECT 280.040 50.225 280.330 50.270 ;
        RECT 283.160 50.225 283.450 50.270 ;
        RECT 285.050 50.225 285.340 50.270 ;
        RECT 280.040 50.085 285.340 50.225 ;
        RECT 280.040 50.040 280.330 50.085 ;
        RECT 283.160 50.040 283.450 50.085 ;
        RECT 285.050 50.040 285.340 50.085 ;
        RECT 303.815 50.225 304.105 50.270 ;
        RECT 306.595 50.225 306.885 50.270 ;
        RECT 308.455 50.225 308.745 50.270 ;
        RECT 303.815 50.085 308.745 50.225 ;
        RECT 303.815 50.040 304.105 50.085 ;
        RECT 306.595 50.040 306.885 50.085 ;
        RECT 308.455 50.040 308.745 50.085 ;
        RECT 271.645 49.885 271.965 49.945 ;
        RECT 275.325 49.885 275.645 49.945 ;
        RECT 268.055 49.745 275.645 49.885 ;
        RECT 249.565 49.685 249.885 49.745 ;
        RECT 250.960 49.700 251.250 49.745 ;
        RECT 260.145 49.685 260.465 49.745 ;
        RECT 271.645 49.685 271.965 49.745 ;
        RECT 275.325 49.685 275.645 49.745 ;
        RECT 277.180 49.885 277.470 49.930 ;
        RECT 279.465 49.885 279.785 49.945 ;
        RECT 309.825 49.885 310.145 49.945 ;
        RECT 277.180 49.745 310.145 49.885 ;
        RECT 277.180 49.700 277.470 49.745 ;
        RECT 279.465 49.685 279.785 49.745 ;
        RECT 309.825 49.685 310.145 49.745 ;
        RECT 162.095 49.065 311.135 49.545 ;
        RECT 175.520 48.865 175.810 48.910 ;
        RECT 176.425 48.865 176.745 48.925 ;
        RECT 175.520 48.725 176.745 48.865 ;
        RECT 175.520 48.680 175.810 48.725 ;
        RECT 176.425 48.665 176.745 48.725 ;
        RECT 185.180 48.865 185.470 48.910 ;
        RECT 185.625 48.865 185.945 48.925 ;
        RECT 185.180 48.725 185.945 48.865 ;
        RECT 185.180 48.680 185.470 48.725 ;
        RECT 185.625 48.665 185.945 48.725 ;
        RECT 188.860 48.865 189.150 48.910 ;
        RECT 190.685 48.865 191.005 48.925 ;
        RECT 223.805 48.865 224.125 48.925 ;
        RECT 188.860 48.725 191.005 48.865 ;
        RECT 188.860 48.680 189.150 48.725 ;
        RECT 190.685 48.665 191.005 48.725 ;
        RECT 216.075 48.725 224.125 48.865 ;
        RECT 179.645 48.525 179.965 48.585 ;
        RECT 207.705 48.525 208.025 48.585 ;
        RECT 179.645 48.385 208.025 48.525 ;
        RECT 179.645 48.325 179.965 48.385 ;
        RECT 207.705 48.325 208.025 48.385 ;
        RECT 176.885 48.185 177.205 48.245 ;
        RECT 178.280 48.185 178.570 48.230 ;
        RECT 176.885 48.045 178.570 48.185 ;
        RECT 176.885 47.985 177.205 48.045 ;
        RECT 178.280 48.000 178.570 48.045 ;
        RECT 182.880 48.185 183.170 48.230 ;
        RECT 183.325 48.185 183.645 48.245 ;
        RECT 195.760 48.185 196.050 48.230 ;
        RECT 200.805 48.185 201.125 48.245 ;
        RECT 182.880 48.045 183.645 48.185 ;
        RECT 182.880 48.000 183.170 48.045 ;
        RECT 183.325 47.985 183.645 48.045 ;
        RECT 184.335 48.045 188.615 48.185 ;
        RECT 184.335 47.905 184.475 48.045 ;
        RECT 175.965 47.845 176.285 47.905 ;
        RECT 177.820 47.845 178.110 47.890 ;
        RECT 182.405 47.845 182.725 47.905 ;
        RECT 175.965 47.705 178.110 47.845 ;
        RECT 175.965 47.645 176.285 47.705 ;
        RECT 177.820 47.660 178.110 47.705 ;
        RECT 180.195 47.705 182.725 47.845 ;
        RECT 177.360 47.505 177.650 47.550 ;
        RECT 180.195 47.505 180.335 47.705 ;
        RECT 182.405 47.645 182.725 47.705 ;
        RECT 184.245 47.645 184.565 47.905 ;
        RECT 188.475 47.890 188.615 48.045 ;
        RECT 195.760 48.045 201.125 48.185 ;
        RECT 195.760 48.000 196.050 48.045 ;
        RECT 200.805 47.985 201.125 48.045 ;
        RECT 185.180 47.660 185.470 47.890 ;
        RECT 188.400 47.660 188.690 47.890 ;
        RECT 198.505 47.845 198.825 47.905 ;
        RECT 199.440 47.845 199.730 47.890 ;
        RECT 198.505 47.705 199.730 47.845 ;
        RECT 173.065 47.365 180.335 47.505 ;
        RECT 180.565 47.505 180.885 47.565 ;
        RECT 181.960 47.505 182.250 47.550 ;
        RECT 184.705 47.505 185.025 47.565 ;
        RECT 185.255 47.505 185.395 47.660 ;
        RECT 198.505 47.645 198.825 47.705 ;
        RECT 199.440 47.660 199.730 47.705 ;
        RECT 214.145 47.645 214.465 47.905 ;
        RECT 215.080 47.845 215.370 47.890 ;
        RECT 215.525 47.845 215.845 47.905 ;
        RECT 216.075 47.890 216.215 48.725 ;
        RECT 223.805 48.665 224.125 48.725 ;
        RECT 225.185 48.665 225.505 48.925 ;
        RECT 231.625 48.665 231.945 48.925 ;
        RECT 240.840 48.865 241.130 48.910 ;
        RECT 242.205 48.865 242.525 48.925 ;
        RECT 247.725 48.865 248.045 48.925 ;
        RECT 254.625 48.865 254.945 48.925 ;
        RECT 240.840 48.725 242.525 48.865 ;
        RECT 240.840 48.680 241.130 48.725 ;
        RECT 242.205 48.665 242.525 48.725 ;
        RECT 242.755 48.725 254.945 48.865 ;
        RECT 217.330 48.525 217.620 48.570 ;
        RECT 219.220 48.525 219.510 48.570 ;
        RECT 222.340 48.525 222.630 48.570 ;
        RECT 217.330 48.385 222.630 48.525 ;
        RECT 217.330 48.340 217.620 48.385 ;
        RECT 219.220 48.340 219.510 48.385 ;
        RECT 222.340 48.340 222.630 48.385 ;
        RECT 232.970 48.525 233.260 48.570 ;
        RECT 234.860 48.525 235.150 48.570 ;
        RECT 237.980 48.525 238.270 48.570 ;
        RECT 232.970 48.385 238.270 48.525 ;
        RECT 232.970 48.340 233.260 48.385 ;
        RECT 234.860 48.340 235.150 48.385 ;
        RECT 237.980 48.340 238.270 48.385 ;
        RECT 241.285 48.525 241.605 48.585 ;
        RECT 242.755 48.525 242.895 48.725 ;
        RECT 247.725 48.665 248.045 48.725 ;
        RECT 254.625 48.665 254.945 48.725 ;
        RECT 264.760 48.865 265.050 48.910 ;
        RECT 266.140 48.865 266.430 48.910 ;
        RECT 266.585 48.865 266.905 48.925 ;
        RECT 264.760 48.725 266.905 48.865 ;
        RECT 264.760 48.680 265.050 48.725 ;
        RECT 266.140 48.680 266.430 48.725 ;
        RECT 266.585 48.665 266.905 48.725 ;
        RECT 267.060 48.865 267.350 48.910 ;
        RECT 267.505 48.865 267.825 48.925 ;
        RECT 267.060 48.725 267.825 48.865 ;
        RECT 267.060 48.680 267.350 48.725 ;
        RECT 267.505 48.665 267.825 48.725 ;
        RECT 282.240 48.865 282.530 48.910 ;
        RECT 286.825 48.865 287.145 48.925 ;
        RECT 282.240 48.725 287.145 48.865 ;
        RECT 282.240 48.680 282.530 48.725 ;
        RECT 286.825 48.665 287.145 48.725 ;
        RECT 241.285 48.385 242.895 48.525 ;
        RECT 244.160 48.525 244.450 48.570 ;
        RECT 247.280 48.525 247.570 48.570 ;
        RECT 249.170 48.525 249.460 48.570 ;
        RECT 244.160 48.385 249.460 48.525 ;
        RECT 241.285 48.325 241.605 48.385 ;
        RECT 244.160 48.340 244.450 48.385 ;
        RECT 247.280 48.340 247.570 48.385 ;
        RECT 249.170 48.340 249.460 48.385 ;
        RECT 256.890 48.525 257.180 48.570 ;
        RECT 258.780 48.525 259.070 48.570 ;
        RECT 261.900 48.525 262.190 48.570 ;
        RECT 271.200 48.525 271.490 48.570 ;
        RECT 256.890 48.385 262.190 48.525 ;
        RECT 256.890 48.340 257.180 48.385 ;
        RECT 258.780 48.340 259.070 48.385 ;
        RECT 261.900 48.340 262.190 48.385 ;
        RECT 262.535 48.385 271.490 48.525 ;
        RECT 216.460 48.185 216.750 48.230 ;
        RECT 223.805 48.185 224.125 48.245 ;
        RECT 227.485 48.185 227.805 48.245 ;
        RECT 216.460 48.045 227.805 48.185 ;
        RECT 216.460 48.000 216.750 48.045 ;
        RECT 215.080 47.705 215.845 47.845 ;
        RECT 215.080 47.660 215.370 47.705 ;
        RECT 215.525 47.645 215.845 47.705 ;
        RECT 216.000 47.660 216.290 47.890 ;
        RECT 180.565 47.365 182.250 47.505 ;
        RECT 172.285 47.165 172.605 47.225 ;
        RECT 173.065 47.165 173.205 47.365 ;
        RECT 177.360 47.320 177.650 47.365 ;
        RECT 180.565 47.305 180.885 47.365 ;
        RECT 181.960 47.320 182.250 47.365 ;
        RECT 182.955 47.365 185.395 47.505 ;
        RECT 214.235 47.505 214.375 47.645 ;
        RECT 216.535 47.505 216.675 48.000 ;
        RECT 223.805 47.985 224.125 48.045 ;
        RECT 227.485 47.985 227.805 48.045 ;
        RECT 227.945 48.185 228.265 48.245 ;
        RECT 232.100 48.185 232.390 48.230 ;
        RECT 227.945 48.045 232.390 48.185 ;
        RECT 227.945 47.985 228.265 48.045 ;
        RECT 232.100 48.000 232.390 48.045 ;
        RECT 233.480 48.185 233.770 48.230 ;
        RECT 239.905 48.185 240.225 48.245 ;
        RECT 233.480 48.045 240.225 48.185 ;
        RECT 233.480 48.000 233.770 48.045 ;
        RECT 239.905 47.985 240.225 48.045 ;
        RECT 260.145 48.185 260.465 48.245 ;
        RECT 262.535 48.185 262.675 48.385 ;
        RECT 271.200 48.340 271.490 48.385 ;
        RECT 284.490 48.525 284.780 48.570 ;
        RECT 286.380 48.525 286.670 48.570 ;
        RECT 289.500 48.525 289.790 48.570 ;
        RECT 284.490 48.385 289.790 48.525 ;
        RECT 284.490 48.340 284.780 48.385 ;
        RECT 286.380 48.340 286.670 48.385 ;
        RECT 289.500 48.340 289.790 48.385 ;
        RECT 260.145 48.045 262.675 48.185 ;
        RECT 264.285 48.185 264.605 48.245 ;
        RECT 267.505 48.185 267.825 48.245 ;
        RECT 271.275 48.185 271.415 48.340 ;
        RECT 290.505 48.325 290.825 48.585 ;
        RECT 279.020 48.185 279.310 48.230 ;
        RECT 264.285 48.045 267.825 48.185 ;
        RECT 260.145 47.985 260.465 48.045 ;
        RECT 264.285 47.985 264.605 48.045 ;
        RECT 267.505 47.985 267.825 48.045 ;
        RECT 269.895 48.045 270.955 48.185 ;
        RECT 271.275 48.045 279.310 48.185 ;
        RECT 216.925 47.845 217.215 47.890 ;
        RECT 218.760 47.845 219.050 47.890 ;
        RECT 222.340 47.845 222.630 47.890 ;
        RECT 216.925 47.705 222.630 47.845 ;
        RECT 216.925 47.660 217.215 47.705 ;
        RECT 218.760 47.660 219.050 47.705 ;
        RECT 222.340 47.660 222.630 47.705 ;
        RECT 223.420 47.550 223.710 47.865 ;
        RECT 228.865 47.645 229.185 47.905 ;
        RECT 232.565 47.845 232.855 47.890 ;
        RECT 234.400 47.845 234.690 47.890 ;
        RECT 237.980 47.845 238.270 47.890 ;
        RECT 243.125 47.865 243.445 47.905 ;
        RECT 232.565 47.705 238.270 47.845 ;
        RECT 232.565 47.660 232.855 47.705 ;
        RECT 234.400 47.660 234.690 47.705 ;
        RECT 237.980 47.660 238.270 47.705 ;
        RECT 239.060 47.845 239.350 47.865 ;
        RECT 243.080 47.845 243.445 47.865 ;
        RECT 239.060 47.705 243.445 47.845 ;
        RECT 214.235 47.365 216.675 47.505 ;
        RECT 182.955 47.225 183.095 47.365 ;
        RECT 184.705 47.305 185.025 47.365 ;
        RECT 217.840 47.320 218.130 47.550 ;
        RECT 220.120 47.505 220.770 47.550 ;
        RECT 223.420 47.505 224.010 47.550 ;
        RECT 226.105 47.505 226.425 47.565 ;
        RECT 229.325 47.505 229.645 47.565 ;
        RECT 239.060 47.550 239.350 47.705 ;
        RECT 243.080 47.645 243.445 47.705 ;
        RECT 244.160 47.845 244.450 47.890 ;
        RECT 247.740 47.845 248.030 47.890 ;
        RECT 249.575 47.845 249.865 47.890 ;
        RECT 244.160 47.705 249.865 47.845 ;
        RECT 244.160 47.660 244.450 47.705 ;
        RECT 247.740 47.660 248.030 47.705 ;
        RECT 249.575 47.660 249.865 47.705 ;
        RECT 250.025 47.845 250.345 47.905 ;
        RECT 252.800 47.845 253.090 47.890 ;
        RECT 255.545 47.845 255.865 47.905 ;
        RECT 256.020 47.845 256.310 47.890 ;
        RECT 250.025 47.705 256.310 47.845 ;
        RECT 250.025 47.645 250.345 47.705 ;
        RECT 252.800 47.660 253.090 47.705 ;
        RECT 255.545 47.645 255.865 47.705 ;
        RECT 256.020 47.660 256.310 47.705 ;
        RECT 256.485 47.845 256.775 47.890 ;
        RECT 258.320 47.845 258.610 47.890 ;
        RECT 261.900 47.845 262.190 47.890 ;
        RECT 256.485 47.705 262.190 47.845 ;
        RECT 256.485 47.660 256.775 47.705 ;
        RECT 258.320 47.660 258.610 47.705 ;
        RECT 261.900 47.660 262.190 47.705 ;
        RECT 243.080 47.550 243.370 47.645 ;
        RECT 220.120 47.365 229.645 47.505 ;
        RECT 220.120 47.320 220.770 47.365 ;
        RECT 223.720 47.320 224.010 47.365 ;
        RECT 172.285 47.025 173.205 47.165 ;
        RECT 179.185 47.165 179.505 47.225 ;
        RECT 179.660 47.165 179.950 47.210 ;
        RECT 179.185 47.025 179.950 47.165 ;
        RECT 172.285 46.965 172.605 47.025 ;
        RECT 179.185 46.965 179.505 47.025 ;
        RECT 179.660 46.980 179.950 47.025 ;
        RECT 181.500 47.165 181.790 47.210 ;
        RECT 182.865 47.165 183.185 47.225 ;
        RECT 181.500 47.025 183.185 47.165 ;
        RECT 181.500 46.980 181.790 47.025 ;
        RECT 182.865 46.965 183.185 47.025 ;
        RECT 214.160 47.165 214.450 47.210 ;
        RECT 217.365 47.165 217.685 47.225 ;
        RECT 214.160 47.025 217.685 47.165 ;
        RECT 217.915 47.165 218.055 47.320 ;
        RECT 226.105 47.305 226.425 47.365 ;
        RECT 229.325 47.305 229.645 47.365 ;
        RECT 235.760 47.505 236.410 47.550 ;
        RECT 239.060 47.505 239.650 47.550 ;
        RECT 235.760 47.365 239.650 47.505 ;
        RECT 235.760 47.320 236.410 47.365 ;
        RECT 239.360 47.320 239.650 47.365 ;
        RECT 242.780 47.505 243.370 47.550 ;
        RECT 246.020 47.505 246.670 47.550 ;
        RECT 242.780 47.365 246.670 47.505 ;
        RECT 242.780 47.320 243.070 47.365 ;
        RECT 246.020 47.320 246.670 47.365 ;
        RECT 248.645 47.305 248.965 47.565 ;
        RECT 257.385 47.305 257.705 47.565 ;
        RECT 262.980 47.550 263.270 47.865 ;
        RECT 269.360 47.845 269.650 47.890 ;
        RECT 269.895 47.845 270.035 48.045 ;
        RECT 268.055 47.705 270.035 47.845 ;
        RECT 259.680 47.505 260.330 47.550 ;
        RECT 262.980 47.505 263.570 47.550 ;
        RECT 257.935 47.365 263.570 47.505 ;
        RECT 222.425 47.165 222.745 47.225 ;
        RECT 217.915 47.025 222.745 47.165 ;
        RECT 214.160 46.980 214.450 47.025 ;
        RECT 217.365 46.965 217.685 47.025 ;
        RECT 222.425 46.965 222.745 47.025 ;
        RECT 241.300 47.165 241.590 47.210 ;
        RECT 244.965 47.165 245.285 47.225 ;
        RECT 241.300 47.025 245.285 47.165 ;
        RECT 241.300 46.980 241.590 47.025 ;
        RECT 244.965 46.965 245.285 47.025 ;
        RECT 251.865 47.165 252.185 47.225 ;
        RECT 255.545 47.165 255.865 47.225 ;
        RECT 257.935 47.165 258.075 47.365 ;
        RECT 259.680 47.320 260.330 47.365 ;
        RECT 263.280 47.320 263.570 47.365 ;
        RECT 265.205 47.305 265.525 47.565 ;
        RECT 266.300 47.505 266.590 47.550 ;
        RECT 268.055 47.505 268.195 47.705 ;
        RECT 269.360 47.660 269.650 47.705 ;
        RECT 270.280 47.660 270.570 47.890 ;
        RECT 270.815 47.845 270.955 48.045 ;
        RECT 279.020 48.000 279.310 48.045 ;
        RECT 279.465 48.185 279.785 48.245 ;
        RECT 279.940 48.185 280.230 48.230 ;
        RECT 279.465 48.045 280.230 48.185 ;
        RECT 279.465 47.985 279.785 48.045 ;
        RECT 279.940 48.000 280.230 48.045 ;
        RECT 283.620 48.185 283.910 48.230 ;
        RECT 290.595 48.185 290.735 48.325 ;
        RECT 283.620 48.045 290.735 48.185 ;
        RECT 292.360 48.185 292.650 48.230 ;
        RECT 295.580 48.185 295.870 48.230 ;
        RECT 292.360 48.045 295.870 48.185 ;
        RECT 283.620 48.000 283.910 48.045 ;
        RECT 292.360 48.000 292.650 48.045 ;
        RECT 295.580 48.000 295.870 48.045 ;
        RECT 271.660 47.845 271.950 47.890 ;
        RECT 273.025 47.845 273.345 47.905 ;
        RECT 270.815 47.705 273.345 47.845 ;
        RECT 271.660 47.660 271.950 47.705 ;
        RECT 266.300 47.365 268.195 47.505 ;
        RECT 268.440 47.505 268.730 47.550 ;
        RECT 268.885 47.505 269.205 47.565 ;
        RECT 268.440 47.365 269.205 47.505 ;
        RECT 266.300 47.320 266.590 47.365 ;
        RECT 268.440 47.320 268.730 47.365 ;
        RECT 268.885 47.305 269.205 47.365 ;
        RECT 251.865 47.025 258.075 47.165 ;
        RECT 265.295 47.165 265.435 47.305 ;
        RECT 270.355 47.165 270.495 47.660 ;
        RECT 273.025 47.645 273.345 47.705 ;
        RECT 280.385 47.645 280.705 47.905 ;
        RECT 284.085 47.845 284.375 47.890 ;
        RECT 285.920 47.845 286.210 47.890 ;
        RECT 289.500 47.845 289.790 47.890 ;
        RECT 284.085 47.705 289.790 47.845 ;
        RECT 284.085 47.660 284.375 47.705 ;
        RECT 285.920 47.660 286.210 47.705 ;
        RECT 289.500 47.660 289.790 47.705 ;
        RECT 290.580 47.550 290.870 47.865 ;
        RECT 285.000 47.320 285.290 47.550 ;
        RECT 287.280 47.505 287.930 47.550 ;
        RECT 290.580 47.505 291.170 47.550 ;
        RECT 291.425 47.505 291.745 47.565 ;
        RECT 294.185 47.505 294.505 47.565 ;
        RECT 287.280 47.365 294.505 47.505 ;
        RECT 287.280 47.320 287.930 47.365 ;
        RECT 290.880 47.320 291.170 47.365 ;
        RECT 265.295 47.025 270.495 47.165 ;
        RECT 285.075 47.165 285.215 47.320 ;
        RECT 291.425 47.305 291.745 47.365 ;
        RECT 294.185 47.305 294.505 47.365 ;
        RECT 291.885 47.165 292.205 47.225 ;
        RECT 285.075 47.025 292.205 47.165 ;
        RECT 251.865 46.965 252.185 47.025 ;
        RECT 255.545 46.965 255.865 47.025 ;
        RECT 291.885 46.965 292.205 47.025 ;
        RECT 292.805 46.965 293.125 47.225 ;
        RECT 162.095 46.345 311.135 46.825 ;
        RECT 175.045 46.145 175.365 46.205 ;
        RECT 173.065 46.005 175.365 46.145 ;
        RECT 173.065 45.805 173.205 46.005 ;
        RECT 175.045 45.945 175.365 46.005 ;
        RECT 181.500 46.145 181.790 46.190 ;
        RECT 182.865 46.145 183.185 46.205 ;
        RECT 181.500 46.005 183.185 46.145 ;
        RECT 181.500 45.960 181.790 46.005 ;
        RECT 182.865 45.945 183.185 46.005 ;
        RECT 198.965 45.945 199.285 46.205 ;
        RECT 217.825 46.145 218.145 46.205 ;
        RECT 218.300 46.145 218.590 46.190 ;
        RECT 217.825 46.005 218.590 46.145 ;
        RECT 217.825 45.945 218.145 46.005 ;
        RECT 218.300 45.960 218.590 46.005 ;
        RECT 222.885 46.145 223.205 46.205 ;
        RECT 243.125 46.145 243.445 46.205 ;
        RECT 222.885 46.005 241.975 46.145 ;
        RECT 222.885 45.945 223.205 46.005 ;
        RECT 172.835 45.665 173.205 45.805 ;
        RECT 176.420 45.805 177.070 45.850 ;
        RECT 180.020 45.805 180.310 45.850 ;
        RECT 176.420 45.665 180.310 45.805 ;
        RECT 165.845 45.125 166.165 45.185 ;
        RECT 172.835 45.170 172.975 45.665 ;
        RECT 176.420 45.620 177.070 45.665 ;
        RECT 179.720 45.620 180.310 45.665 ;
        RECT 193.900 45.805 194.550 45.850 ;
        RECT 197.500 45.805 197.790 45.850 ;
        RECT 198.045 45.805 198.365 45.865 ;
        RECT 193.900 45.665 198.365 45.805 ;
        RECT 193.900 45.620 194.550 45.665 ;
        RECT 197.200 45.620 197.790 45.665 ;
        RECT 173.225 45.465 173.515 45.510 ;
        RECT 175.060 45.465 175.350 45.510 ;
        RECT 178.640 45.465 178.930 45.510 ;
        RECT 173.225 45.325 178.930 45.465 ;
        RECT 173.225 45.280 173.515 45.325 ;
        RECT 175.060 45.280 175.350 45.325 ;
        RECT 178.640 45.280 178.930 45.325 ;
        RECT 179.720 45.465 180.010 45.620 ;
        RECT 183.785 45.465 184.105 45.525 ;
        RECT 179.720 45.325 184.105 45.465 ;
        RECT 179.720 45.305 180.010 45.325 ;
        RECT 183.785 45.265 184.105 45.325 ;
        RECT 189.305 45.265 189.625 45.525 ;
        RECT 190.705 45.465 190.995 45.510 ;
        RECT 192.540 45.465 192.830 45.510 ;
        RECT 196.120 45.465 196.410 45.510 ;
        RECT 190.705 45.325 196.410 45.465 ;
        RECT 190.705 45.280 190.995 45.325 ;
        RECT 192.540 45.280 192.830 45.325 ;
        RECT 196.120 45.280 196.410 45.325 ;
        RECT 197.200 45.305 197.490 45.620 ;
        RECT 198.045 45.605 198.365 45.665 ;
        RECT 209.545 45.805 209.865 45.865 ;
        RECT 229.785 45.805 230.105 45.865 ;
        RECT 209.545 45.665 230.105 45.805 ;
        RECT 209.545 45.605 209.865 45.665 ;
        RECT 198.965 45.465 199.285 45.525 ;
        RECT 200.820 45.465 201.110 45.510 ;
        RECT 198.965 45.325 201.110 45.465 ;
        RECT 198.965 45.265 199.285 45.325 ;
        RECT 200.820 45.280 201.110 45.325 ;
        RECT 204.485 45.465 204.805 45.525 ;
        RECT 204.485 45.325 217.595 45.465 ;
        RECT 204.485 45.265 204.805 45.325 ;
        RECT 172.760 45.125 173.050 45.170 ;
        RECT 165.845 44.985 173.050 45.125 ;
        RECT 165.845 44.925 166.165 44.985 ;
        RECT 172.760 44.940 173.050 44.985 ;
        RECT 174.140 45.125 174.430 45.170 ;
        RECT 179.185 45.125 179.505 45.185 ;
        RECT 174.140 44.985 179.505 45.125 ;
        RECT 174.140 44.940 174.430 44.985 ;
        RECT 179.185 44.925 179.505 44.985 ;
        RECT 180.565 45.125 180.885 45.185 ;
        RECT 182.420 45.125 182.710 45.170 ;
        RECT 180.565 44.985 182.710 45.125 ;
        RECT 180.565 44.925 180.885 44.985 ;
        RECT 182.420 44.940 182.710 44.985 ;
        RECT 185.165 44.925 185.485 45.185 ;
        RECT 190.240 44.940 190.530 45.170 ;
        RECT 191.620 45.125 191.910 45.170 ;
        RECT 207.705 45.125 208.025 45.185 ;
        RECT 212.765 45.125 213.085 45.185 ;
        RECT 191.620 44.985 203.335 45.125 ;
        RECT 191.620 44.940 191.910 44.985 ;
        RECT 173.630 44.785 173.920 44.830 ;
        RECT 175.520 44.785 175.810 44.830 ;
        RECT 178.640 44.785 178.930 44.830 ;
        RECT 187.465 44.785 187.785 44.845 ;
        RECT 190.315 44.785 190.455 44.940 ;
        RECT 173.630 44.645 178.930 44.785 ;
        RECT 173.630 44.600 173.920 44.645 ;
        RECT 175.520 44.600 175.810 44.645 ;
        RECT 178.640 44.600 178.930 44.645 ;
        RECT 181.115 44.645 190.455 44.785 ;
        RECT 175.045 44.445 175.365 44.505 ;
        RECT 181.115 44.445 181.255 44.645 ;
        RECT 187.465 44.585 187.785 44.645 ;
        RECT 175.045 44.305 181.255 44.445 ;
        RECT 185.625 44.445 185.945 44.505 ;
        RECT 187.925 44.445 188.245 44.505 ;
        RECT 188.860 44.445 189.150 44.490 ;
        RECT 185.625 44.305 189.150 44.445 ;
        RECT 190.315 44.445 190.455 44.645 ;
        RECT 191.110 44.785 191.400 44.830 ;
        RECT 193.000 44.785 193.290 44.830 ;
        RECT 196.120 44.785 196.410 44.830 ;
        RECT 191.110 44.645 196.410 44.785 ;
        RECT 191.110 44.600 191.400 44.645 ;
        RECT 193.000 44.600 193.290 44.645 ;
        RECT 196.120 44.600 196.410 44.645 ;
        RECT 202.645 44.585 202.965 44.845 ;
        RECT 193.905 44.445 194.225 44.505 ;
        RECT 203.195 44.490 203.335 44.985 ;
        RECT 207.705 44.985 217.135 45.125 ;
        RECT 207.705 44.925 208.025 44.985 ;
        RECT 212.765 44.925 213.085 44.985 ;
        RECT 190.315 44.305 194.225 44.445 ;
        RECT 175.045 44.245 175.365 44.305 ;
        RECT 185.625 44.245 185.945 44.305 ;
        RECT 187.925 44.245 188.245 44.305 ;
        RECT 188.860 44.260 189.150 44.305 ;
        RECT 193.905 44.245 194.225 44.305 ;
        RECT 203.120 44.445 203.410 44.490 ;
        RECT 207.245 44.445 207.565 44.505 ;
        RECT 203.120 44.305 207.565 44.445 ;
        RECT 203.120 44.260 203.410 44.305 ;
        RECT 207.245 44.245 207.565 44.305 ;
        RECT 216.445 44.245 216.765 44.505 ;
        RECT 216.995 44.445 217.135 44.985 ;
        RECT 217.455 44.785 217.595 45.325 ;
        RECT 218.745 44.925 219.065 45.185 ;
        RECT 219.295 45.170 219.435 45.665 ;
        RECT 229.785 45.605 230.105 45.665 ;
        RECT 233.920 45.805 234.570 45.850 ;
        RECT 237.520 45.805 237.810 45.850 ;
        RECT 233.920 45.665 237.810 45.805 ;
        RECT 233.920 45.620 234.570 45.665 ;
        RECT 237.220 45.620 237.810 45.665 ;
        RECT 237.220 45.525 237.510 45.620 ;
        RECT 223.805 45.265 224.125 45.525 ;
        RECT 224.725 45.265 225.045 45.525 ;
        RECT 225.185 45.465 225.505 45.525 ;
        RECT 227.500 45.465 227.790 45.510 ;
        RECT 225.185 45.325 227.790 45.465 ;
        RECT 225.185 45.265 225.505 45.325 ;
        RECT 227.500 45.280 227.790 45.325 ;
        RECT 228.405 45.265 228.725 45.525 ;
        RECT 230.260 45.280 230.550 45.510 ;
        RECT 230.725 45.465 231.015 45.510 ;
        RECT 232.560 45.465 232.850 45.510 ;
        RECT 236.140 45.465 236.430 45.510 ;
        RECT 230.725 45.325 236.430 45.465 ;
        RECT 230.725 45.280 231.015 45.325 ;
        RECT 232.560 45.280 232.850 45.325 ;
        RECT 236.140 45.280 236.430 45.325 ;
        RECT 237.145 45.305 237.510 45.525 ;
        RECT 240.840 45.465 241.130 45.510 ;
        RECT 241.285 45.465 241.605 45.525 ;
        RECT 241.835 45.510 241.975 46.005 ;
        RECT 243.125 46.005 251.175 46.145 ;
        RECT 243.125 45.945 243.445 46.005 ;
        RECT 242.205 45.805 242.525 45.865 ;
        RECT 250.025 45.805 250.345 45.865 ;
        RECT 242.205 45.665 247.035 45.805 ;
        RECT 242.205 45.605 242.525 45.665 ;
        RECT 237.695 45.325 241.605 45.465 ;
        RECT 219.220 44.940 219.510 45.170 ;
        RECT 223.345 44.785 223.665 44.845 ;
        RECT 217.455 44.645 223.665 44.785 ;
        RECT 223.345 44.585 223.665 44.645 ;
        RECT 223.805 44.785 224.125 44.845 ;
        RECT 227.945 44.785 228.265 44.845 ;
        RECT 230.335 44.785 230.475 45.280 ;
        RECT 237.145 45.265 237.465 45.305 ;
        RECT 231.640 45.125 231.930 45.170 ;
        RECT 232.085 45.125 232.405 45.185 ;
        RECT 231.640 44.985 232.405 45.125 ;
        RECT 231.640 44.940 231.930 44.985 ;
        RECT 232.085 44.925 232.405 44.985 ;
        RECT 235.305 45.125 235.625 45.185 ;
        RECT 237.695 45.125 237.835 45.325 ;
        RECT 240.840 45.280 241.130 45.325 ;
        RECT 241.285 45.265 241.605 45.325 ;
        RECT 241.760 45.280 242.050 45.510 ;
        RECT 242.665 45.265 242.985 45.525 ;
        RECT 243.600 45.465 243.890 45.510 ;
        RECT 246.345 45.465 246.665 45.525 ;
        RECT 246.895 45.510 247.035 45.665 ;
        RECT 248.275 45.665 250.345 45.805 ;
        RECT 251.035 45.805 251.175 46.005 ;
        RECT 257.385 45.945 257.705 46.205 ;
        RECT 268.440 46.145 268.730 46.190 ;
        RECT 265.295 46.005 268.730 46.145 ;
        RECT 265.295 45.865 265.435 46.005 ;
        RECT 268.440 45.960 268.730 46.005 ;
        RECT 273.025 45.945 273.345 46.205 ;
        RECT 280.385 46.145 280.705 46.205 ;
        RECT 282.240 46.145 282.530 46.190 ;
        RECT 280.385 46.005 282.530 46.145 ;
        RECT 280.385 45.945 280.705 46.005 ;
        RECT 282.240 45.960 282.530 46.005 ;
        RECT 251.865 45.850 252.185 45.865 ;
        RECT 251.860 45.805 252.510 45.850 ;
        RECT 255.460 45.805 255.750 45.850 ;
        RECT 265.205 45.805 265.525 45.865 ;
        RECT 251.035 45.665 255.750 45.805 ;
        RECT 248.275 45.510 248.415 45.665 ;
        RECT 250.025 45.605 250.345 45.665 ;
        RECT 251.860 45.620 252.510 45.665 ;
        RECT 255.160 45.620 255.750 45.665 ;
        RECT 258.855 45.665 265.525 45.805 ;
        RECT 251.865 45.605 252.185 45.620 ;
        RECT 243.600 45.325 246.665 45.465 ;
        RECT 243.600 45.280 243.890 45.325 ;
        RECT 246.345 45.265 246.665 45.325 ;
        RECT 246.820 45.280 247.110 45.510 ;
        RECT 248.200 45.280 248.490 45.510 ;
        RECT 248.665 45.465 248.955 45.510 ;
        RECT 250.500 45.465 250.790 45.510 ;
        RECT 254.080 45.465 254.370 45.510 ;
        RECT 248.665 45.325 254.370 45.465 ;
        RECT 248.665 45.280 248.955 45.325 ;
        RECT 250.500 45.280 250.790 45.325 ;
        RECT 254.080 45.280 254.370 45.325 ;
        RECT 255.160 45.305 255.450 45.620 ;
        RECT 258.320 45.465 258.610 45.510 ;
        RECT 258.855 45.465 258.995 45.665 ;
        RECT 265.205 45.605 265.525 45.665 ;
        RECT 266.585 45.605 266.905 45.865 ;
        RECT 267.505 45.605 267.825 45.865 ;
        RECT 300.160 45.805 300.810 45.850 ;
        RECT 303.760 45.805 304.050 45.850 ;
        RECT 300.160 45.665 304.050 45.805 ;
        RECT 300.160 45.620 300.810 45.665 ;
        RECT 303.460 45.620 304.050 45.665 ;
        RECT 258.320 45.325 258.995 45.465 ;
        RECT 258.320 45.280 258.610 45.325 ;
        RECT 235.305 44.985 237.835 45.125 ;
        RECT 235.305 44.925 235.625 44.985 ;
        RECT 238.985 44.925 239.305 45.185 ;
        RECT 242.220 45.125 242.510 45.170 ;
        RECT 244.060 45.125 244.350 45.170 ;
        RECT 242.220 44.985 244.350 45.125 ;
        RECT 242.220 44.940 242.510 44.985 ;
        RECT 244.060 44.940 244.350 44.985 ;
        RECT 249.565 44.925 249.885 45.185 ;
        RECT 254.625 45.125 254.945 45.185 ;
        RECT 258.395 45.125 258.535 45.280 ;
        RECT 259.225 45.265 259.545 45.525 ;
        RECT 260.145 45.265 260.465 45.525 ;
        RECT 261.080 45.465 261.370 45.510 ;
        RECT 265.680 45.465 265.970 45.510 ;
        RECT 261.080 45.325 265.970 45.465 ;
        RECT 261.080 45.280 261.370 45.325 ;
        RECT 265.680 45.280 265.970 45.325 ;
        RECT 267.980 45.465 268.270 45.510 ;
        RECT 268.885 45.465 269.205 45.525 ;
        RECT 267.980 45.325 269.205 45.465 ;
        RECT 267.980 45.280 268.270 45.325 ;
        RECT 268.885 45.265 269.205 45.325 ;
        RECT 271.660 45.465 271.950 45.510 ;
        RECT 272.105 45.465 272.425 45.525 ;
        RECT 271.660 45.325 272.425 45.465 ;
        RECT 271.660 45.280 271.950 45.325 ;
        RECT 272.105 45.265 272.425 45.325 ;
        RECT 272.655 45.325 275.095 45.465 ;
        RECT 254.625 44.985 258.535 45.125 ;
        RECT 259.700 45.125 259.990 45.170 ;
        RECT 261.540 45.125 261.830 45.170 ;
        RECT 259.700 44.985 261.830 45.125 ;
        RECT 254.625 44.925 254.945 44.985 ;
        RECT 259.700 44.940 259.990 44.985 ;
        RECT 261.540 44.940 261.830 44.985 ;
        RECT 264.300 44.940 264.590 45.170 ;
        RECT 269.805 45.125 270.125 45.185 ;
        RECT 272.655 45.125 272.795 45.325 ;
        RECT 269.805 44.985 272.795 45.125 ;
        RECT 273.040 45.125 273.330 45.170 ;
        RECT 274.405 45.125 274.725 45.185 ;
        RECT 273.040 44.985 274.725 45.125 ;
        RECT 223.805 44.645 230.475 44.785 ;
        RECT 231.130 44.785 231.420 44.830 ;
        RECT 233.020 44.785 233.310 44.830 ;
        RECT 236.140 44.785 236.430 44.830 ;
        RECT 231.130 44.645 236.430 44.785 ;
        RECT 223.805 44.585 224.125 44.645 ;
        RECT 227.945 44.585 228.265 44.645 ;
        RECT 231.130 44.600 231.420 44.645 ;
        RECT 233.020 44.600 233.310 44.645 ;
        RECT 236.140 44.600 236.430 44.645 ;
        RECT 239.920 44.785 240.210 44.830 ;
        RECT 244.505 44.785 244.825 44.845 ;
        RECT 239.920 44.645 244.825 44.785 ;
        RECT 239.920 44.600 240.210 44.645 ;
        RECT 244.505 44.585 244.825 44.645 ;
        RECT 249.070 44.785 249.360 44.830 ;
        RECT 250.960 44.785 251.250 44.830 ;
        RECT 254.080 44.785 254.370 44.830 ;
        RECT 249.070 44.645 254.370 44.785 ;
        RECT 249.070 44.600 249.360 44.645 ;
        RECT 250.960 44.600 251.250 44.645 ;
        RECT 254.080 44.600 254.370 44.645 ;
        RECT 256.925 44.785 257.245 44.845 ;
        RECT 264.375 44.785 264.515 44.940 ;
        RECT 269.805 44.925 270.125 44.985 ;
        RECT 273.040 44.940 273.330 44.985 ;
        RECT 274.405 44.925 274.725 44.985 ;
        RECT 256.925 44.645 264.515 44.785 ;
        RECT 264.745 44.785 265.065 44.845 ;
        RECT 273.960 44.785 274.250 44.830 ;
        RECT 264.745 44.645 274.250 44.785 ;
        RECT 256.925 44.585 257.245 44.645 ;
        RECT 264.745 44.585 265.065 44.645 ;
        RECT 273.960 44.600 274.250 44.645 ;
        RECT 228.405 44.445 228.725 44.505 ;
        RECT 216.995 44.305 228.725 44.445 ;
        RECT 228.405 44.245 228.725 44.305 ;
        RECT 229.325 44.445 229.645 44.505 ;
        RECT 232.545 44.445 232.865 44.505 ;
        RECT 229.325 44.305 232.865 44.445 ;
        RECT 229.325 44.245 229.645 44.305 ;
        RECT 232.545 44.245 232.865 44.305 ;
        RECT 255.545 44.445 255.865 44.505 ;
        RECT 267.505 44.445 267.825 44.505 ;
        RECT 255.545 44.305 267.825 44.445 ;
        RECT 255.545 44.245 255.865 44.305 ;
        RECT 267.505 44.245 267.825 44.305 ;
        RECT 270.725 44.445 271.045 44.505 ;
        RECT 272.120 44.445 272.410 44.490 ;
        RECT 270.725 44.305 272.410 44.445 ;
        RECT 274.955 44.445 275.095 45.325 ;
        RECT 279.005 45.265 279.325 45.525 ;
        RECT 296.965 45.465 297.255 45.510 ;
        RECT 298.800 45.465 299.090 45.510 ;
        RECT 302.380 45.465 302.670 45.510 ;
        RECT 296.965 45.325 302.670 45.465 ;
        RECT 296.965 45.280 297.255 45.325 ;
        RECT 298.800 45.280 299.090 45.325 ;
        RECT 302.380 45.280 302.670 45.325 ;
        RECT 303.460 45.465 303.750 45.620 ;
        RECT 304.305 45.465 304.625 45.525 ;
        RECT 303.460 45.325 304.625 45.465 ;
        RECT 303.460 45.305 303.750 45.325 ;
        RECT 304.305 45.265 304.625 45.325 ;
        RECT 305.225 45.465 305.545 45.525 ;
        RECT 308.000 45.465 308.290 45.510 ;
        RECT 305.225 45.325 308.290 45.465 ;
        RECT 305.225 45.265 305.545 45.325 ;
        RECT 308.000 45.280 308.290 45.325 ;
        RECT 277.180 45.125 277.470 45.170 ;
        RECT 285.445 45.125 285.765 45.185 ;
        RECT 277.180 44.985 285.765 45.125 ;
        RECT 277.180 44.940 277.470 44.985 ;
        RECT 285.445 44.925 285.765 44.985 ;
        RECT 285.905 45.125 286.225 45.185 ;
        RECT 296.485 45.125 296.805 45.185 ;
        RECT 285.905 44.985 296.805 45.125 ;
        RECT 285.905 44.925 286.225 44.985 ;
        RECT 296.485 44.925 296.805 44.985 ;
        RECT 297.880 45.125 298.170 45.170 ;
        RECT 310.285 45.125 310.605 45.185 ;
        RECT 297.880 44.985 310.605 45.125 ;
        RECT 297.880 44.940 298.170 44.985 ;
        RECT 310.285 44.925 310.605 44.985 ;
        RECT 297.370 44.785 297.660 44.830 ;
        RECT 299.260 44.785 299.550 44.830 ;
        RECT 302.380 44.785 302.670 44.830 ;
        RECT 297.370 44.645 302.670 44.785 ;
        RECT 297.370 44.600 297.660 44.645 ;
        RECT 299.260 44.600 299.550 44.645 ;
        RECT 302.380 44.600 302.670 44.645 ;
        RECT 304.305 44.785 304.625 44.845 ;
        RECT 308.920 44.785 309.210 44.830 ;
        RECT 304.305 44.645 309.210 44.785 ;
        RECT 304.305 44.585 304.625 44.645 ;
        RECT 308.920 44.600 309.210 44.645 ;
        RECT 304.765 44.445 305.085 44.505 ;
        RECT 274.955 44.305 305.085 44.445 ;
        RECT 270.725 44.245 271.045 44.305 ;
        RECT 272.120 44.260 272.410 44.305 ;
        RECT 304.765 44.245 305.085 44.305 ;
        RECT 305.240 44.445 305.530 44.490 ;
        RECT 306.145 44.445 306.465 44.505 ;
        RECT 305.240 44.305 306.465 44.445 ;
        RECT 305.240 44.260 305.530 44.305 ;
        RECT 306.145 44.245 306.465 44.305 ;
        RECT 162.095 43.625 311.135 44.105 ;
        RECT 174.600 43.425 174.890 43.470 ;
        RECT 185.165 43.425 185.485 43.485 ;
        RECT 174.600 43.285 185.485 43.425 ;
        RECT 174.600 43.240 174.890 43.285 ;
        RECT 185.165 43.225 185.485 43.285 ;
        RECT 210.005 43.425 210.325 43.485 ;
        RECT 223.820 43.425 224.110 43.470 ;
        RECT 224.265 43.425 224.585 43.485 ;
        RECT 210.005 43.285 213.455 43.425 ;
        RECT 210.005 43.225 210.325 43.285 ;
        RECT 166.730 43.085 167.020 43.130 ;
        RECT 168.620 43.085 168.910 43.130 ;
        RECT 171.740 43.085 172.030 43.130 ;
        RECT 166.730 42.945 172.030 43.085 ;
        RECT 166.730 42.900 167.020 42.945 ;
        RECT 168.620 42.900 168.910 42.945 ;
        RECT 171.740 42.900 172.030 42.945 ;
        RECT 176.390 43.085 176.680 43.130 ;
        RECT 178.280 43.085 178.570 43.130 ;
        RECT 181.400 43.085 181.690 43.130 ;
        RECT 176.390 42.945 181.690 43.085 ;
        RECT 176.390 42.900 176.680 42.945 ;
        RECT 178.280 42.900 178.570 42.945 ;
        RECT 181.400 42.900 181.690 42.945 ;
        RECT 189.880 43.085 190.170 43.130 ;
        RECT 193.000 43.085 193.290 43.130 ;
        RECT 194.890 43.085 195.180 43.130 ;
        RECT 189.880 42.945 195.180 43.085 ;
        RECT 189.880 42.900 190.170 42.945 ;
        RECT 193.000 42.900 193.290 42.945 ;
        RECT 194.890 42.900 195.180 42.945 ;
        RECT 202.150 43.085 202.440 43.130 ;
        RECT 204.040 43.085 204.330 43.130 ;
        RECT 207.160 43.085 207.450 43.130 ;
        RECT 202.150 42.945 207.450 43.085 ;
        RECT 202.150 42.900 202.440 42.945 ;
        RECT 204.040 42.900 204.330 42.945 ;
        RECT 207.160 42.900 207.450 42.945 ;
        RECT 175.045 42.745 175.365 42.805 ;
        RECT 175.520 42.745 175.810 42.790 ;
        RECT 175.045 42.605 175.810 42.745 ;
        RECT 175.045 42.545 175.365 42.605 ;
        RECT 175.520 42.560 175.810 42.605 ;
        RECT 195.760 42.745 196.050 42.790 ;
        RECT 200.805 42.745 201.125 42.805 ;
        RECT 213.315 42.790 213.455 43.285 ;
        RECT 223.820 43.285 224.585 43.425 ;
        RECT 223.820 43.240 224.110 43.285 ;
        RECT 224.265 43.225 224.585 43.285 ;
        RECT 228.865 43.425 229.185 43.485 ;
        RECT 234.860 43.425 235.150 43.470 ;
        RECT 228.865 43.285 235.150 43.425 ;
        RECT 228.865 43.225 229.185 43.285 ;
        RECT 234.860 43.240 235.150 43.285 ;
        RECT 247.740 43.425 248.030 43.470 ;
        RECT 248.645 43.425 248.965 43.485 ;
        RECT 247.740 43.285 248.965 43.425 ;
        RECT 247.740 43.240 248.030 43.285 ;
        RECT 248.645 43.225 248.965 43.285 ;
        RECT 256.005 43.225 256.325 43.485 ;
        RECT 269.805 43.425 270.125 43.485 ;
        RECT 256.555 43.285 270.125 43.425 ;
        RECT 215.950 43.085 216.240 43.130 ;
        RECT 217.840 43.085 218.130 43.130 ;
        RECT 220.960 43.085 221.250 43.130 ;
        RECT 215.950 42.945 221.250 43.085 ;
        RECT 215.950 42.900 216.240 42.945 ;
        RECT 217.840 42.900 218.130 42.945 ;
        RECT 220.960 42.900 221.250 42.945 ;
        RECT 223.345 43.085 223.665 43.145 ;
        RECT 240.380 43.085 240.670 43.130 ;
        RECT 242.665 43.085 242.985 43.145 ;
        RECT 245.885 43.085 246.205 43.145 ;
        RECT 223.345 42.945 236.915 43.085 ;
        RECT 223.345 42.885 223.665 42.945 ;
        RECT 201.280 42.745 201.570 42.790 ;
        RECT 195.760 42.605 201.570 42.745 ;
        RECT 195.760 42.560 196.050 42.605 ;
        RECT 200.805 42.545 201.125 42.605 ;
        RECT 201.280 42.560 201.570 42.605 ;
        RECT 213.240 42.560 213.530 42.790 ;
        RECT 214.145 42.745 214.465 42.805 ;
        RECT 215.080 42.745 215.370 42.790 ;
        RECT 223.805 42.745 224.125 42.805 ;
        RECT 236.225 42.745 236.545 42.805 ;
        RECT 236.775 42.790 236.915 42.945 ;
        RECT 240.380 42.945 242.985 43.085 ;
        RECT 240.380 42.900 240.670 42.945 ;
        RECT 242.665 42.885 242.985 42.945 ;
        RECT 243.675 42.945 246.205 43.085 ;
        RECT 214.145 42.605 224.125 42.745 ;
        RECT 214.145 42.545 214.465 42.605 ;
        RECT 215.080 42.560 215.370 42.605 ;
        RECT 223.805 42.545 224.125 42.605 ;
        RECT 224.355 42.605 236.545 42.745 ;
        RECT 165.845 42.205 166.165 42.465 ;
        RECT 166.325 42.405 166.615 42.450 ;
        RECT 168.160 42.405 168.450 42.450 ;
        RECT 171.740 42.405 172.030 42.450 ;
        RECT 166.325 42.265 172.030 42.405 ;
        RECT 166.325 42.220 166.615 42.265 ;
        RECT 168.160 42.220 168.450 42.265 ;
        RECT 171.740 42.220 172.030 42.265 ;
        RECT 172.745 42.425 173.065 42.465 ;
        RECT 172.745 42.205 173.110 42.425 ;
        RECT 175.985 42.405 176.275 42.450 ;
        RECT 177.820 42.405 178.110 42.450 ;
        RECT 181.400 42.405 181.690 42.450 ;
        RECT 175.985 42.265 181.690 42.405 ;
        RECT 175.985 42.220 176.275 42.265 ;
        RECT 177.820 42.220 178.110 42.265 ;
        RECT 181.400 42.220 181.690 42.265 ;
        RECT 172.820 42.110 173.110 42.205 ;
        RECT 167.240 41.880 167.530 42.110 ;
        RECT 169.520 42.065 170.170 42.110 ;
        RECT 172.820 42.065 173.410 42.110 ;
        RECT 169.520 41.925 173.410 42.065 ;
        RECT 169.520 41.880 170.170 41.925 ;
        RECT 173.120 41.880 173.410 41.925 ;
        RECT 176.900 42.065 177.190 42.110 ;
        RECT 177.345 42.065 177.665 42.125 ;
        RECT 182.480 42.110 182.770 42.425 ;
        RECT 176.900 41.925 177.665 42.065 ;
        RECT 176.900 41.880 177.190 41.925 ;
        RECT 167.315 41.725 167.455 41.880 ;
        RECT 177.345 41.865 177.665 41.925 ;
        RECT 179.180 42.065 179.830 42.110 ;
        RECT 182.480 42.065 183.070 42.110 ;
        RECT 183.785 42.065 184.105 42.125 ;
        RECT 188.800 42.110 189.090 42.425 ;
        RECT 189.880 42.405 190.170 42.450 ;
        RECT 193.460 42.405 193.750 42.450 ;
        RECT 195.295 42.405 195.585 42.450 ;
        RECT 189.880 42.265 195.585 42.405 ;
        RECT 189.880 42.220 190.170 42.265 ;
        RECT 193.460 42.220 193.750 42.265 ;
        RECT 195.295 42.220 195.585 42.265 ;
        RECT 201.745 42.405 202.035 42.450 ;
        RECT 203.580 42.405 203.870 42.450 ;
        RECT 207.160 42.405 207.450 42.450 ;
        RECT 201.745 42.265 207.450 42.405 ;
        RECT 201.745 42.220 202.035 42.265 ;
        RECT 203.580 42.220 203.870 42.265 ;
        RECT 207.160 42.220 207.450 42.265 ;
        RECT 179.180 41.925 184.105 42.065 ;
        RECT 179.180 41.880 179.830 41.925 ;
        RECT 182.780 41.880 183.070 41.925 ;
        RECT 183.785 41.865 184.105 41.925 ;
        RECT 188.500 42.065 189.090 42.110 ;
        RECT 191.740 42.065 192.390 42.110 ;
        RECT 192.985 42.065 193.305 42.125 ;
        RECT 188.500 41.925 194.135 42.065 ;
        RECT 188.500 41.880 188.790 41.925 ;
        RECT 191.740 41.880 192.390 41.925 ;
        RECT 192.985 41.865 193.305 41.925 ;
        RECT 175.505 41.725 175.825 41.785 ;
        RECT 167.315 41.585 175.825 41.725 ;
        RECT 175.505 41.525 175.825 41.585 ;
        RECT 184.245 41.525 184.565 41.785 ;
        RECT 187.005 41.525 187.325 41.785 ;
        RECT 193.995 41.725 194.135 41.925 ;
        RECT 194.365 41.865 194.685 42.125 ;
        RECT 202.660 42.065 202.950 42.110 ;
        RECT 204.025 42.065 204.345 42.125 ;
        RECT 208.240 42.110 208.530 42.425 ;
        RECT 215.545 42.405 215.835 42.450 ;
        RECT 217.380 42.405 217.670 42.450 ;
        RECT 220.960 42.405 221.250 42.450 ;
        RECT 215.545 42.265 221.250 42.405 ;
        RECT 215.545 42.220 215.835 42.265 ;
        RECT 217.380 42.220 217.670 42.265 ;
        RECT 220.960 42.220 221.250 42.265 ;
        RECT 221.965 42.425 222.285 42.465 ;
        RECT 221.965 42.405 222.330 42.425 ;
        RECT 224.355 42.405 224.495 42.605 ;
        RECT 236.225 42.545 236.545 42.605 ;
        RECT 236.700 42.560 236.990 42.790 ;
        RECT 242.205 42.745 242.525 42.805 ;
        RECT 243.675 42.790 243.815 42.945 ;
        RECT 245.885 42.885 246.205 42.945 ;
        RECT 246.345 43.085 246.665 43.145 ;
        RECT 248.200 43.085 248.490 43.130 ;
        RECT 256.555 43.085 256.695 43.285 ;
        RECT 269.805 43.225 270.125 43.285 ;
        RECT 274.405 43.225 274.725 43.485 ;
        RECT 246.345 42.945 248.490 43.085 ;
        RECT 246.345 42.885 246.665 42.945 ;
        RECT 248.200 42.900 248.490 42.945 ;
        RECT 249.655 42.945 256.695 43.085 ;
        RECT 266.550 43.085 266.840 43.130 ;
        RECT 268.440 43.085 268.730 43.130 ;
        RECT 271.560 43.085 271.850 43.130 ;
        RECT 266.550 42.945 271.850 43.085 ;
        RECT 237.695 42.605 242.525 42.745 ;
        RECT 221.965 42.265 224.495 42.405 ;
        RECT 224.725 42.405 225.045 42.465 ;
        RECT 228.880 42.405 229.170 42.450 ;
        RECT 224.725 42.265 229.170 42.405 ;
        RECT 221.965 42.205 222.330 42.265 ;
        RECT 224.725 42.205 225.045 42.265 ;
        RECT 228.880 42.220 229.170 42.265 ;
        RECT 233.465 42.205 233.785 42.465 ;
        RECT 235.305 42.405 235.625 42.465 ;
        RECT 235.780 42.405 236.070 42.450 ;
        RECT 235.305 42.265 236.070 42.405 ;
        RECT 235.305 42.205 235.625 42.265 ;
        RECT 235.780 42.220 236.070 42.265 ;
        RECT 237.145 42.205 237.465 42.465 ;
        RECT 237.695 42.450 237.835 42.605 ;
        RECT 242.205 42.545 242.525 42.605 ;
        RECT 243.600 42.560 243.890 42.790 ;
        RECT 244.505 42.545 244.825 42.805 ;
        RECT 237.620 42.220 237.910 42.450 ;
        RECT 238.540 42.220 238.830 42.450 ;
        RECT 244.965 42.405 245.285 42.465 ;
        RECT 249.120 42.405 249.410 42.450 ;
        RECT 244.965 42.265 249.410 42.405 ;
        RECT 202.660 41.925 204.345 42.065 ;
        RECT 202.660 41.880 202.950 41.925 ;
        RECT 204.025 41.865 204.345 41.925 ;
        RECT 204.940 42.065 205.590 42.110 ;
        RECT 208.240 42.065 208.830 42.110 ;
        RECT 209.085 42.065 209.405 42.125 ;
        RECT 204.940 41.925 209.405 42.065 ;
        RECT 204.940 41.880 205.590 41.925 ;
        RECT 208.540 41.880 208.830 41.925 ;
        RECT 209.085 41.865 209.405 41.925 ;
        RECT 216.445 41.865 216.765 42.125 ;
        RECT 222.040 42.110 222.330 42.205 ;
        RECT 218.740 42.065 219.390 42.110 ;
        RECT 222.040 42.065 222.630 42.110 ;
        RECT 227.040 42.065 227.330 42.110 ;
        RECT 238.615 42.065 238.755 42.220 ;
        RECT 244.965 42.205 245.285 42.265 ;
        RECT 249.120 42.220 249.410 42.265 ;
        RECT 218.740 41.925 222.630 42.065 ;
        RECT 218.740 41.880 219.390 41.925 ;
        RECT 222.340 41.880 222.630 41.925 ;
        RECT 223.435 41.925 227.330 42.065 ;
        RECT 198.045 41.725 198.365 41.785 ;
        RECT 193.995 41.585 198.365 41.725 ;
        RECT 198.045 41.525 198.365 41.585 ;
        RECT 210.465 41.525 210.785 41.785 ;
        RECT 217.825 41.725 218.145 41.785 ;
        RECT 223.435 41.725 223.575 41.925 ;
        RECT 227.040 41.880 227.330 41.925 ;
        RECT 229.415 41.925 238.755 42.065 ;
        RECT 241.835 41.925 243.815 42.065 ;
        RECT 217.825 41.585 223.575 41.725 ;
        RECT 226.565 41.725 226.885 41.785 ;
        RECT 229.415 41.725 229.555 41.925 ;
        RECT 226.565 41.585 229.555 41.725 ;
        RECT 230.720 41.725 231.010 41.770 ;
        RECT 232.085 41.725 232.405 41.785 ;
        RECT 230.720 41.585 232.405 41.725 ;
        RECT 217.825 41.525 218.145 41.585 ;
        RECT 226.565 41.525 226.885 41.585 ;
        RECT 230.720 41.540 231.010 41.585 ;
        RECT 232.085 41.525 232.405 41.585 ;
        RECT 238.525 41.725 238.845 41.785 ;
        RECT 241.835 41.725 241.975 41.925 ;
        RECT 238.525 41.585 241.975 41.725 ;
        RECT 238.525 41.525 238.845 41.585 ;
        RECT 242.205 41.525 242.525 41.785 ;
        RECT 242.680 41.725 242.970 41.770 ;
        RECT 243.125 41.725 243.445 41.785 ;
        RECT 242.680 41.585 243.445 41.725 ;
        RECT 243.675 41.725 243.815 41.925 ;
        RECT 249.655 41.725 249.795 42.945 ;
        RECT 266.550 42.900 266.840 42.945 ;
        RECT 268.440 42.900 268.730 42.945 ;
        RECT 271.560 42.900 271.850 42.945 ;
        RECT 288.320 43.085 288.610 43.130 ;
        RECT 291.440 43.085 291.730 43.130 ;
        RECT 293.330 43.085 293.620 43.130 ;
        RECT 288.320 42.945 293.620 43.085 ;
        RECT 288.320 42.900 288.610 42.945 ;
        RECT 291.440 42.900 291.730 42.945 ;
        RECT 293.330 42.900 293.620 42.945 ;
        RECT 265.680 42.745 265.970 42.790 ;
        RECT 258.855 42.605 265.970 42.745 ;
        RECT 258.855 42.465 258.995 42.605 ;
        RECT 265.680 42.560 265.970 42.605 ;
        RECT 267.505 42.745 267.825 42.805 ;
        RECT 267.505 42.605 273.255 42.745 ;
        RECT 267.505 42.545 267.825 42.605 ;
        RECT 250.040 42.405 250.330 42.450 ;
        RECT 250.945 42.405 251.265 42.465 ;
        RECT 250.040 42.265 251.265 42.405 ;
        RECT 250.040 42.220 250.330 42.265 ;
        RECT 250.945 42.205 251.265 42.265 ;
        RECT 255.100 42.405 255.390 42.450 ;
        RECT 256.005 42.405 256.325 42.465 ;
        RECT 258.765 42.405 259.085 42.465 ;
        RECT 255.100 42.265 259.085 42.405 ;
        RECT 255.100 42.220 255.390 42.265 ;
        RECT 256.005 42.205 256.325 42.265 ;
        RECT 258.765 42.205 259.085 42.265 ;
        RECT 259.225 42.205 259.545 42.465 ;
        RECT 260.160 42.405 260.450 42.450 ;
        RECT 262.905 42.405 263.225 42.465 ;
        RECT 260.160 42.265 263.225 42.405 ;
        RECT 260.160 42.220 260.450 42.265 ;
        RECT 262.905 42.205 263.225 42.265 ;
        RECT 266.145 42.405 266.435 42.450 ;
        RECT 267.980 42.405 268.270 42.450 ;
        RECT 271.560 42.405 271.850 42.450 ;
        RECT 266.145 42.265 271.850 42.405 ;
        RECT 266.145 42.220 266.435 42.265 ;
        RECT 267.980 42.220 268.270 42.265 ;
        RECT 271.560 42.220 271.850 42.265 ;
        RECT 243.675 41.585 249.795 41.725 ;
        RECT 251.035 41.725 251.175 42.205 ;
        RECT 256.925 41.865 257.245 42.125 ;
        RECT 257.860 42.065 258.150 42.110 ;
        RECT 264.285 42.065 264.605 42.125 ;
        RECT 257.860 41.925 264.605 42.065 ;
        RECT 257.860 41.880 258.150 41.925 ;
        RECT 257.935 41.725 258.075 41.880 ;
        RECT 264.285 41.865 264.605 41.925 ;
        RECT 265.205 42.065 265.525 42.125 ;
        RECT 272.640 42.110 272.930 42.425 ;
        RECT 273.115 42.110 273.255 42.605 ;
        RECT 285.460 42.560 285.750 42.790 ;
        RECT 290.505 42.745 290.825 42.805 ;
        RECT 294.200 42.745 294.490 42.790 ;
        RECT 290.505 42.605 294.490 42.745 ;
        RECT 281.305 42.405 281.625 42.465 ;
        RECT 285.535 42.405 285.675 42.560 ;
        RECT 290.505 42.545 290.825 42.605 ;
        RECT 294.200 42.560 294.490 42.605 ;
        RECT 306.145 42.545 306.465 42.805 ;
        RECT 281.305 42.265 285.675 42.405 ;
        RECT 281.305 42.205 281.625 42.265 ;
        RECT 267.060 42.065 267.350 42.110 ;
        RECT 265.205 41.925 267.350 42.065 ;
        RECT 265.205 41.865 265.525 41.925 ;
        RECT 267.060 41.880 267.350 41.925 ;
        RECT 269.340 42.065 269.990 42.110 ;
        RECT 272.640 42.065 273.255 42.110 ;
        RECT 274.880 42.065 275.170 42.110 ;
        RECT 269.340 41.925 275.170 42.065 ;
        RECT 269.340 41.880 269.990 41.925 ;
        RECT 272.940 41.880 273.230 41.925 ;
        RECT 274.880 41.880 275.170 41.925 ;
        RECT 276.705 42.065 277.025 42.125 ;
        RECT 287.240 42.110 287.530 42.425 ;
        RECT 288.320 42.405 288.610 42.450 ;
        RECT 291.900 42.405 292.190 42.450 ;
        RECT 293.735 42.405 294.025 42.450 ;
        RECT 288.320 42.265 294.025 42.405 ;
        RECT 288.320 42.220 288.610 42.265 ;
        RECT 291.900 42.220 292.190 42.265 ;
        RECT 293.735 42.220 294.025 42.265 ;
        RECT 304.765 42.405 305.085 42.465 ;
        RECT 307.065 42.405 307.385 42.465 ;
        RECT 304.765 42.265 307.385 42.405 ;
        RECT 304.765 42.205 305.085 42.265 ;
        RECT 307.065 42.205 307.385 42.265 ;
        RECT 286.940 42.065 287.530 42.110 ;
        RECT 290.180 42.065 290.830 42.110 ;
        RECT 291.425 42.065 291.745 42.125 ;
        RECT 276.705 41.925 279.235 42.065 ;
        RECT 276.705 41.865 277.025 41.925 ;
        RECT 251.035 41.585 258.075 41.725 ;
        RECT 258.305 41.725 258.625 41.785 ;
        RECT 259.700 41.725 259.990 41.770 ;
        RECT 258.305 41.585 259.990 41.725 ;
        RECT 242.680 41.540 242.970 41.585 ;
        RECT 243.125 41.525 243.445 41.585 ;
        RECT 258.305 41.525 258.625 41.585 ;
        RECT 259.700 41.540 259.990 41.585 ;
        RECT 270.725 41.725 271.045 41.785 ;
        RECT 277.625 41.725 277.945 41.785 ;
        RECT 270.725 41.585 277.945 41.725 ;
        RECT 270.725 41.525 271.045 41.585 ;
        RECT 277.625 41.525 277.945 41.585 ;
        RECT 278.085 41.725 278.405 41.785 ;
        RECT 278.560 41.725 278.850 41.770 ;
        RECT 278.085 41.585 278.850 41.725 ;
        RECT 279.095 41.725 279.235 41.925 ;
        RECT 286.940 41.925 291.745 42.065 ;
        RECT 286.940 41.880 287.230 41.925 ;
        RECT 290.180 41.880 290.830 41.925 ;
        RECT 291.425 41.865 291.745 41.925 ;
        RECT 292.805 41.865 293.125 42.125 ;
        RECT 305.225 41.725 305.545 41.785 ;
        RECT 279.095 41.585 305.545 41.725 ;
        RECT 278.085 41.525 278.405 41.585 ;
        RECT 278.560 41.540 278.850 41.585 ;
        RECT 305.225 41.525 305.545 41.585 ;
        RECT 307.065 41.725 307.385 41.785 ;
        RECT 309.380 41.725 309.670 41.770 ;
        RECT 307.065 41.585 309.670 41.725 ;
        RECT 307.065 41.525 307.385 41.585 ;
        RECT 309.380 41.540 309.670 41.585 ;
        RECT 162.095 40.905 311.135 41.385 ;
        RECT 177.345 40.505 177.665 40.765 ;
        RECT 179.200 40.705 179.490 40.750 ;
        RECT 184.245 40.705 184.565 40.765 ;
        RECT 179.200 40.565 184.565 40.705 ;
        RECT 179.200 40.520 179.490 40.565 ;
        RECT 184.245 40.505 184.565 40.565 ;
        RECT 185.625 40.505 185.945 40.765 ;
        RECT 189.780 40.705 190.070 40.750 ;
        RECT 194.365 40.705 194.685 40.765 ;
        RECT 200.805 40.705 201.125 40.765 ;
        RECT 189.780 40.565 194.685 40.705 ;
        RECT 189.780 40.520 190.070 40.565 ;
        RECT 194.365 40.505 194.685 40.565 ;
        RECT 195.375 40.565 201.125 40.705 ;
        RECT 171.820 40.365 172.470 40.410 ;
        RECT 175.420 40.365 175.710 40.410 ;
        RECT 183.785 40.365 184.105 40.425 ;
        RECT 171.820 40.225 184.105 40.365 ;
        RECT 171.820 40.180 172.470 40.225 ;
        RECT 175.120 40.180 175.735 40.225 ;
        RECT 168.625 40.025 168.915 40.070 ;
        RECT 170.460 40.025 170.750 40.070 ;
        RECT 174.040 40.025 174.330 40.070 ;
        RECT 168.625 39.885 174.330 40.025 ;
        RECT 168.625 39.840 168.915 39.885 ;
        RECT 170.460 39.840 170.750 39.885 ;
        RECT 174.040 39.840 174.330 39.885 ;
        RECT 175.120 39.865 175.410 40.180 ;
        RECT 167.685 39.685 168.005 39.745 ;
        RECT 168.160 39.685 168.450 39.730 ;
        RECT 167.685 39.545 168.450 39.685 ;
        RECT 167.685 39.485 168.005 39.545 ;
        RECT 168.160 39.500 168.450 39.545 ;
        RECT 168.235 39.005 168.375 39.500 ;
        RECT 169.525 39.485 169.845 39.745 ;
        RECT 172.745 39.685 173.065 39.745 ;
        RECT 175.595 39.685 175.735 40.180 ;
        RECT 183.785 40.165 184.105 40.225 ;
        RECT 187.005 40.365 187.325 40.425 ;
        RECT 191.620 40.365 191.910 40.410 ;
        RECT 187.005 40.225 191.910 40.365 ;
        RECT 187.005 40.165 187.325 40.225 ;
        RECT 191.620 40.180 191.910 40.225 ;
        RECT 195.375 40.070 195.515 40.565 ;
        RECT 200.805 40.505 201.125 40.565 ;
        RECT 204.025 40.705 204.345 40.765 ;
        RECT 204.500 40.705 204.790 40.750 ;
        RECT 204.025 40.565 204.790 40.705 ;
        RECT 204.025 40.505 204.345 40.565 ;
        RECT 204.500 40.520 204.790 40.565 ;
        RECT 206.340 40.705 206.630 40.750 ;
        RECT 210.465 40.705 210.785 40.765 ;
        RECT 206.340 40.565 210.785 40.705 ;
        RECT 206.340 40.520 206.630 40.565 ;
        RECT 210.465 40.505 210.785 40.565 ;
        RECT 217.365 40.705 217.685 40.765 ;
        RECT 226.565 40.705 226.885 40.765 ;
        RECT 217.365 40.565 226.885 40.705 ;
        RECT 217.365 40.505 217.685 40.565 ;
        RECT 226.565 40.505 226.885 40.565 ;
        RECT 227.500 40.705 227.790 40.750 ;
        RECT 232.085 40.705 232.405 40.765 ;
        RECT 227.500 40.565 232.405 40.705 ;
        RECT 227.500 40.520 227.790 40.565 ;
        RECT 232.085 40.505 232.405 40.565 ;
        RECT 237.145 40.505 237.465 40.765 ;
        RECT 242.205 40.705 242.525 40.765 ;
        RECT 247.740 40.705 248.030 40.750 ;
        RECT 264.745 40.705 265.065 40.765 ;
        RECT 272.580 40.705 272.870 40.750 ;
        RECT 242.205 40.565 265.065 40.705 ;
        RECT 242.205 40.505 242.525 40.565 ;
        RECT 247.740 40.520 248.030 40.565 ;
        RECT 264.745 40.505 265.065 40.565 ;
        RECT 269.665 40.565 272.870 40.705 ;
        RECT 198.045 40.365 198.365 40.425 ;
        RECT 198.960 40.365 199.610 40.410 ;
        RECT 202.560 40.365 202.850 40.410 ;
        RECT 198.045 40.225 202.850 40.365 ;
        RECT 198.045 40.165 198.365 40.225 ;
        RECT 198.960 40.180 199.610 40.225 ;
        RECT 202.260 40.180 202.850 40.225 ;
        RECT 217.820 40.365 218.470 40.410 ;
        RECT 221.420 40.365 221.710 40.410 ;
        RECT 221.965 40.365 222.285 40.425 ;
        RECT 217.820 40.225 222.285 40.365 ;
        RECT 217.820 40.180 218.470 40.225 ;
        RECT 221.120 40.180 221.710 40.225 ;
        RECT 195.300 39.840 195.590 40.070 ;
        RECT 195.765 40.025 196.055 40.070 ;
        RECT 197.600 40.025 197.890 40.070 ;
        RECT 201.180 40.025 201.470 40.070 ;
        RECT 195.765 39.885 201.470 40.025 ;
        RECT 195.765 39.840 196.055 39.885 ;
        RECT 197.600 39.840 197.890 39.885 ;
        RECT 201.180 39.840 201.470 39.885 ;
        RECT 202.260 39.865 202.550 40.180 ;
        RECT 206.800 40.025 207.090 40.070 ;
        RECT 208.625 40.025 208.945 40.085 ;
        RECT 206.800 39.885 208.945 40.025 ;
        RECT 206.800 39.840 207.090 39.885 ;
        RECT 208.625 39.825 208.945 39.885 ;
        RECT 214.145 39.825 214.465 40.085 ;
        RECT 214.625 40.025 214.915 40.070 ;
        RECT 216.460 40.025 216.750 40.070 ;
        RECT 220.040 40.025 220.330 40.070 ;
        RECT 214.625 39.885 220.330 40.025 ;
        RECT 214.625 39.840 214.915 39.885 ;
        RECT 216.460 39.840 216.750 39.885 ;
        RECT 220.040 39.840 220.330 39.885 ;
        RECT 221.120 39.865 221.410 40.180 ;
        RECT 221.965 40.165 222.285 40.225 ;
        RECT 222.885 40.365 223.205 40.425 ;
        RECT 224.280 40.365 224.570 40.410 ;
        RECT 222.885 40.225 224.570 40.365 ;
        RECT 222.885 40.165 223.205 40.225 ;
        RECT 224.280 40.180 224.570 40.225 ;
        RECT 225.200 40.365 225.490 40.410 ;
        RECT 225.645 40.365 225.965 40.425 ;
        RECT 225.200 40.225 225.965 40.365 ;
        RECT 225.200 40.180 225.490 40.225 ;
        RECT 225.645 40.165 225.965 40.225 ;
        RECT 228.405 40.365 228.725 40.425 ;
        RECT 237.620 40.365 237.910 40.410 ;
        RECT 243.140 40.365 243.430 40.410 ;
        RECT 245.425 40.365 245.745 40.425 ;
        RECT 228.405 40.225 237.910 40.365 ;
        RECT 228.405 40.165 228.725 40.225 ;
        RECT 237.620 40.180 237.910 40.225 ;
        RECT 238.155 40.225 241.515 40.365 ;
        RECT 231.640 40.025 231.930 40.070 ;
        RECT 233.005 40.025 233.325 40.085 ;
        RECT 238.155 40.025 238.295 40.225 ;
        RECT 231.640 39.885 233.325 40.025 ;
        RECT 231.640 39.840 231.930 39.885 ;
        RECT 233.005 39.825 233.325 39.885 ;
        RECT 234.015 39.885 238.295 40.025 ;
        RECT 172.745 39.545 175.735 39.685 ;
        RECT 175.965 39.685 176.285 39.745 ;
        RECT 179.660 39.685 179.950 39.730 ;
        RECT 175.965 39.545 179.950 39.685 ;
        RECT 172.745 39.485 173.065 39.545 ;
        RECT 175.965 39.485 176.285 39.545 ;
        RECT 179.660 39.500 179.950 39.545 ;
        RECT 180.580 39.685 180.870 39.730 ;
        RECT 183.325 39.685 183.645 39.745 ;
        RECT 180.580 39.545 185.855 39.685 ;
        RECT 180.580 39.500 180.870 39.545 ;
        RECT 183.325 39.485 183.645 39.545 ;
        RECT 169.030 39.345 169.320 39.390 ;
        RECT 170.920 39.345 171.210 39.390 ;
        RECT 174.040 39.345 174.330 39.390 ;
        RECT 184.245 39.345 184.565 39.405 ;
        RECT 169.030 39.205 174.330 39.345 ;
        RECT 169.030 39.160 169.320 39.205 ;
        RECT 170.920 39.160 171.210 39.205 ;
        RECT 174.040 39.160 174.330 39.205 ;
        RECT 176.515 39.205 184.565 39.345 ;
        RECT 185.715 39.345 185.855 39.545 ;
        RECT 186.085 39.485 186.405 39.745 ;
        RECT 187.020 39.500 187.310 39.730 ;
        RECT 187.095 39.345 187.235 39.500 ;
        RECT 192.065 39.485 192.385 39.745 ;
        RECT 193.000 39.685 193.290 39.730 ;
        RECT 196.680 39.685 196.970 39.730 ;
        RECT 198.505 39.685 198.825 39.745 ;
        RECT 193.000 39.545 195.975 39.685 ;
        RECT 193.000 39.500 193.290 39.545 ;
        RECT 193.075 39.345 193.215 39.500 ;
        RECT 185.715 39.205 193.215 39.345 ;
        RECT 176.515 39.005 176.655 39.205 ;
        RECT 184.245 39.145 184.565 39.205 ;
        RECT 168.235 38.865 176.655 39.005 ;
        RECT 176.885 38.805 177.205 39.065 ;
        RECT 183.800 39.005 184.090 39.050 ;
        RECT 185.625 39.005 185.945 39.065 ;
        RECT 183.800 38.865 185.945 39.005 ;
        RECT 195.835 39.005 195.975 39.545 ;
        RECT 196.680 39.545 198.825 39.685 ;
        RECT 196.680 39.500 196.970 39.545 ;
        RECT 198.505 39.485 198.825 39.545 ;
        RECT 202.645 39.685 202.965 39.745 ;
        RECT 204.040 39.685 204.330 39.730 ;
        RECT 202.645 39.545 204.330 39.685 ;
        RECT 202.645 39.485 202.965 39.545 ;
        RECT 204.040 39.500 204.330 39.545 ;
        RECT 207.245 39.685 207.565 39.745 ;
        RECT 209.545 39.685 209.865 39.745 ;
        RECT 207.245 39.545 209.865 39.685 ;
        RECT 207.245 39.485 207.565 39.545 ;
        RECT 209.545 39.485 209.865 39.545 ;
        RECT 210.480 39.500 210.770 39.730 ;
        RECT 213.240 39.685 213.530 39.730 ;
        RECT 215.540 39.685 215.830 39.730 ;
        RECT 213.240 39.545 215.830 39.685 ;
        RECT 213.240 39.500 213.530 39.545 ;
        RECT 215.540 39.500 215.830 39.545 ;
        RECT 218.285 39.685 218.605 39.745 ;
        RECT 223.360 39.685 223.650 39.730 ;
        RECT 218.285 39.545 220.815 39.685 ;
        RECT 196.170 39.345 196.460 39.390 ;
        RECT 198.060 39.345 198.350 39.390 ;
        RECT 201.180 39.345 201.470 39.390 ;
        RECT 196.170 39.205 201.470 39.345 ;
        RECT 196.170 39.160 196.460 39.205 ;
        RECT 198.060 39.160 198.350 39.205 ;
        RECT 201.180 39.160 201.470 39.205 ;
        RECT 207.335 39.005 207.475 39.485 ;
        RECT 195.835 38.865 207.475 39.005 ;
        RECT 210.555 39.005 210.695 39.500 ;
        RECT 218.285 39.485 218.605 39.545 ;
        RECT 215.030 39.345 215.320 39.390 ;
        RECT 216.920 39.345 217.210 39.390 ;
        RECT 220.040 39.345 220.330 39.390 ;
        RECT 215.030 39.205 220.330 39.345 ;
        RECT 220.675 39.345 220.815 39.545 ;
        RECT 222.055 39.545 223.650 39.685 ;
        RECT 222.055 39.345 222.195 39.545 ;
        RECT 223.360 39.500 223.650 39.545 ;
        RECT 227.945 39.485 228.265 39.745 ;
        RECT 228.880 39.500 229.170 39.730 ;
        RECT 229.785 39.685 230.105 39.745 ;
        RECT 232.560 39.685 232.850 39.730 ;
        RECT 234.015 39.685 234.155 39.885 ;
        RECT 238.525 39.825 238.845 40.085 ;
        RECT 229.785 39.545 234.155 39.685 ;
        RECT 234.400 39.685 234.690 39.730 ;
        RECT 238.985 39.685 239.305 39.745 ;
        RECT 234.400 39.545 239.305 39.685 ;
        RECT 241.375 39.685 241.515 40.225 ;
        RECT 243.140 40.225 245.745 40.365 ;
        RECT 243.140 40.180 243.430 40.225 ;
        RECT 245.425 40.165 245.745 40.225 ;
        RECT 254.625 40.165 254.945 40.425 ;
        RECT 255.720 40.365 256.010 40.410 ;
        RECT 262.445 40.365 262.765 40.425 ;
        RECT 268.885 40.365 269.205 40.425 ;
        RECT 255.720 40.225 262.765 40.365 ;
        RECT 255.720 40.180 256.010 40.225 ;
        RECT 262.445 40.165 262.765 40.225 ;
        RECT 265.755 40.225 269.205 40.365 ;
        RECT 243.600 40.025 243.890 40.070 ;
        RECT 247.280 40.025 247.570 40.070 ;
        RECT 249.580 40.025 249.870 40.070 ;
        RECT 256.940 40.025 257.230 40.070 ;
        RECT 243.600 39.885 249.870 40.025 ;
        RECT 243.600 39.840 243.890 39.885 ;
        RECT 247.280 39.840 247.570 39.885 ;
        RECT 249.580 39.840 249.870 39.885 ;
        RECT 250.115 39.885 257.230 40.025 ;
        RECT 244.060 39.685 244.350 39.730 ;
        RECT 241.375 39.545 244.350 39.685 ;
        RECT 228.955 39.345 229.095 39.500 ;
        RECT 229.785 39.485 230.105 39.545 ;
        RECT 232.560 39.500 232.850 39.545 ;
        RECT 234.400 39.500 234.690 39.545 ;
        RECT 238.985 39.485 239.305 39.545 ;
        RECT 244.060 39.500 244.350 39.545 ;
        RECT 248.660 39.685 248.950 39.730 ;
        RECT 250.115 39.685 250.255 39.885 ;
        RECT 256.940 39.840 257.230 39.885 ;
        RECT 258.305 39.825 258.625 40.085 ;
        RECT 258.765 40.025 259.085 40.085 ;
        RECT 260.620 40.025 260.910 40.070 ;
        RECT 258.765 39.885 260.910 40.025 ;
        RECT 258.765 39.825 259.085 39.885 ;
        RECT 260.620 39.840 260.910 39.885 ;
        RECT 248.660 39.545 250.255 39.685 ;
        RECT 248.660 39.500 248.950 39.545 ;
        RECT 248.735 39.345 248.875 39.500 ;
        RECT 252.325 39.485 252.645 39.745 ;
        RECT 260.695 39.685 260.835 39.840 ;
        RECT 261.985 39.825 262.305 40.085 ;
        RECT 265.755 40.025 265.895 40.225 ;
        RECT 268.885 40.165 269.205 40.225 ;
        RECT 269.665 40.025 269.805 40.565 ;
        RECT 272.580 40.520 272.870 40.565 ;
        RECT 273.025 40.705 273.345 40.765 ;
        RECT 278.100 40.705 278.390 40.750 ;
        RECT 281.305 40.705 281.625 40.765 ;
        RECT 273.025 40.565 281.625 40.705 ;
        RECT 273.025 40.505 273.345 40.565 ;
        RECT 278.100 40.520 278.390 40.565 ;
        RECT 281.305 40.505 281.625 40.565 ;
        RECT 296.485 40.705 296.805 40.765 ;
        RECT 296.485 40.565 308.675 40.705 ;
        RECT 296.485 40.505 296.805 40.565 ;
        RECT 304.305 40.410 304.625 40.425 ;
        RECT 301.200 40.365 301.490 40.410 ;
        RECT 304.305 40.365 305.090 40.410 ;
        RECT 262.535 39.885 265.895 40.025 ;
        RECT 266.215 39.885 269.805 40.025 ;
        RECT 270.815 40.225 276.935 40.365 ;
        RECT 262.535 39.685 262.675 39.885 ;
        RECT 252.875 39.545 258.995 39.685 ;
        RECT 260.695 39.545 262.675 39.685 ;
        RECT 263.380 39.685 263.670 39.730 ;
        RECT 265.680 39.685 265.970 39.730 ;
        RECT 263.380 39.545 265.970 39.685 ;
        RECT 220.675 39.205 222.195 39.345 ;
        RECT 222.515 39.205 248.875 39.345 ;
        RECT 215.030 39.160 215.320 39.205 ;
        RECT 216.920 39.160 217.210 39.205 ;
        RECT 220.040 39.160 220.330 39.205 ;
        RECT 214.145 39.005 214.465 39.065 ;
        RECT 210.555 38.865 214.465 39.005 ;
        RECT 183.800 38.820 184.090 38.865 ;
        RECT 185.625 38.805 185.945 38.865 ;
        RECT 214.145 38.805 214.465 38.865 ;
        RECT 221.045 39.005 221.365 39.065 ;
        RECT 222.515 39.005 222.655 39.205 ;
        RECT 221.045 38.865 222.655 39.005 ;
        RECT 221.045 38.805 221.365 38.865 ;
        RECT 222.885 38.805 223.205 39.065 ;
        RECT 225.645 38.805 225.965 39.065 ;
        RECT 229.800 39.005 230.090 39.050 ;
        RECT 230.245 39.005 230.565 39.065 ;
        RECT 229.800 38.865 230.565 39.005 ;
        RECT 229.800 38.820 230.090 38.865 ;
        RECT 230.245 38.805 230.565 38.865 ;
        RECT 241.285 38.805 241.605 39.065 ;
        RECT 242.205 39.005 242.525 39.065 ;
        RECT 245.440 39.005 245.730 39.050 ;
        RECT 242.205 38.865 245.730 39.005 ;
        RECT 242.205 38.805 242.525 38.865 ;
        RECT 245.440 38.820 245.730 38.865 ;
        RECT 245.885 39.005 246.205 39.065 ;
        RECT 252.875 39.005 253.015 39.545 ;
        RECT 258.305 39.345 258.625 39.405 ;
        RECT 255.635 39.205 258.625 39.345 ;
        RECT 258.855 39.345 258.995 39.545 ;
        RECT 263.380 39.500 263.670 39.545 ;
        RECT 265.680 39.500 265.970 39.545 ;
        RECT 266.215 39.345 266.355 39.885 ;
        RECT 267.045 39.685 267.365 39.745 ;
        RECT 268.440 39.685 268.730 39.730 ;
        RECT 270.815 39.685 270.955 40.225 ;
        RECT 271.200 40.025 271.490 40.070 ;
        RECT 276.245 40.025 276.565 40.085 ;
        RECT 271.200 39.885 276.565 40.025 ;
        RECT 271.200 39.840 271.490 39.885 ;
        RECT 267.045 39.545 268.730 39.685 ;
        RECT 267.045 39.485 267.365 39.545 ;
        RECT 268.440 39.500 268.730 39.545 ;
        RECT 269.665 39.545 270.955 39.685 ;
        RECT 271.660 39.685 271.950 39.730 ;
        RECT 272.105 39.685 272.425 39.745 ;
        RECT 274.035 39.730 274.175 39.885 ;
        RECT 276.245 39.825 276.565 39.885 ;
        RECT 271.660 39.545 272.425 39.685 ;
        RECT 269.665 39.345 269.805 39.545 ;
        RECT 271.660 39.500 271.950 39.545 ;
        RECT 272.105 39.485 272.425 39.545 ;
        RECT 273.960 39.500 274.250 39.730 ;
        RECT 274.420 39.685 274.710 39.730 ;
        RECT 274.420 39.545 274.820 39.685 ;
        RECT 274.420 39.500 274.710 39.545 ;
        RECT 275.800 39.500 276.090 39.730 ;
        RECT 274.495 39.345 274.635 39.500 ;
        RECT 275.875 39.345 276.015 39.500 ;
        RECT 276.795 39.390 276.935 40.225 ;
        RECT 301.200 40.225 305.090 40.365 ;
        RECT 301.200 40.180 301.790 40.225 ;
        RECT 277.180 39.840 277.470 40.070 ;
        RECT 277.255 39.685 277.395 39.840 ;
        RECT 277.625 39.825 277.945 40.085 ;
        RECT 279.020 40.025 279.310 40.070 ;
        RECT 279.940 40.025 280.230 40.070 ;
        RECT 279.020 39.885 280.230 40.025 ;
        RECT 279.020 39.840 279.310 39.885 ;
        RECT 279.940 39.840 280.230 39.885 ;
        RECT 301.500 39.865 301.790 40.180 ;
        RECT 304.305 40.180 305.090 40.225 ;
        RECT 304.305 40.165 304.625 40.180 ;
        RECT 307.065 40.165 307.385 40.425 ;
        RECT 308.535 40.070 308.675 40.565 ;
        RECT 302.580 40.025 302.870 40.070 ;
        RECT 306.160 40.025 306.450 40.070 ;
        RECT 307.995 40.025 308.285 40.070 ;
        RECT 302.580 39.885 308.285 40.025 ;
        RECT 302.580 39.840 302.870 39.885 ;
        RECT 306.160 39.840 306.450 39.885 ;
        RECT 307.995 39.840 308.285 39.885 ;
        RECT 308.460 39.840 308.750 40.070 ;
        RECT 277.255 39.545 279.235 39.685 ;
        RECT 279.095 39.390 279.235 39.545 ;
        RECT 282.685 39.485 283.005 39.745 ;
        RECT 285.445 39.685 285.765 39.745 ;
        RECT 299.720 39.685 300.010 39.730 ;
        RECT 285.445 39.545 300.010 39.685 ;
        RECT 285.445 39.485 285.765 39.545 ;
        RECT 299.720 39.500 300.010 39.545 ;
        RECT 258.855 39.205 266.355 39.345 ;
        RECT 266.675 39.205 269.805 39.345 ;
        RECT 270.355 39.205 276.015 39.345 ;
        RECT 255.635 39.050 255.775 39.205 ;
        RECT 258.305 39.145 258.625 39.205 ;
        RECT 266.675 39.065 266.815 39.205 ;
        RECT 245.885 38.865 253.015 39.005 ;
        RECT 245.885 38.805 246.205 38.865 ;
        RECT 255.560 38.820 255.850 39.050 ;
        RECT 256.480 39.005 256.770 39.050 ;
        RECT 256.925 39.005 257.245 39.065 ;
        RECT 256.480 38.865 257.245 39.005 ;
        RECT 256.480 38.820 256.770 38.865 ;
        RECT 256.925 38.805 257.245 38.865 ;
        RECT 257.385 39.005 257.705 39.065 ;
        RECT 261.080 39.005 261.370 39.050 ;
        RECT 257.385 38.865 261.370 39.005 ;
        RECT 257.385 38.805 257.705 38.865 ;
        RECT 261.080 38.820 261.370 38.865 ;
        RECT 262.920 39.005 263.210 39.050 ;
        RECT 266.585 39.005 266.905 39.065 ;
        RECT 262.920 38.865 266.905 39.005 ;
        RECT 262.920 38.820 263.210 38.865 ;
        RECT 266.585 38.805 266.905 38.865 ;
        RECT 268.885 39.005 269.205 39.065 ;
        RECT 270.355 39.005 270.495 39.205 ;
        RECT 276.720 39.160 277.010 39.390 ;
        RECT 279.020 39.160 279.310 39.390 ;
        RECT 302.580 39.345 302.870 39.390 ;
        RECT 305.700 39.345 305.990 39.390 ;
        RECT 307.590 39.345 307.880 39.390 ;
        RECT 302.580 39.205 307.880 39.345 ;
        RECT 302.580 39.160 302.870 39.205 ;
        RECT 305.700 39.160 305.990 39.205 ;
        RECT 307.590 39.160 307.880 39.205 ;
        RECT 268.885 38.865 270.495 39.005 ;
        RECT 268.885 38.805 269.205 38.865 ;
        RECT 270.725 38.805 271.045 39.065 ;
        RECT 273.025 39.005 273.345 39.065 ;
        RECT 276.260 39.005 276.550 39.050 ;
        RECT 273.025 38.865 276.550 39.005 ;
        RECT 276.795 39.005 276.935 39.160 ;
        RECT 281.305 39.005 281.625 39.065 ;
        RECT 276.795 38.865 281.625 39.005 ;
        RECT 273.025 38.805 273.345 38.865 ;
        RECT 276.260 38.820 276.550 38.865 ;
        RECT 281.305 38.805 281.625 38.865 ;
        RECT 283.145 39.005 283.465 39.065 ;
        RECT 291.425 39.005 291.745 39.065 ;
        RECT 283.145 38.865 291.745 39.005 ;
        RECT 283.145 38.805 283.465 38.865 ;
        RECT 291.425 38.805 291.745 38.865 ;
        RECT 162.095 38.185 311.135 38.665 ;
        RECT 167.240 37.985 167.530 38.030 ;
        RECT 169.525 37.985 169.845 38.045 ;
        RECT 167.240 37.845 169.845 37.985 ;
        RECT 167.240 37.800 167.530 37.845 ;
        RECT 169.525 37.785 169.845 37.845 ;
        RECT 175.505 37.785 175.825 38.045 ;
        RECT 183.800 37.985 184.090 38.030 ;
        RECT 186.085 37.985 186.405 38.045 ;
        RECT 183.800 37.845 186.405 37.985 ;
        RECT 183.800 37.800 184.090 37.845 ;
        RECT 186.085 37.785 186.405 37.845 ;
        RECT 189.305 37.985 189.625 38.045 ;
        RECT 193.000 37.985 193.290 38.030 ;
        RECT 189.305 37.845 193.290 37.985 ;
        RECT 189.305 37.785 189.625 37.845 ;
        RECT 193.000 37.800 193.290 37.845 ;
        RECT 214.605 37.985 214.925 38.045 ;
        RECT 215.080 37.985 215.370 38.030 ;
        RECT 214.605 37.845 215.370 37.985 ;
        RECT 214.605 37.785 214.925 37.845 ;
        RECT 215.080 37.800 215.370 37.845 ;
        RECT 218.745 37.985 219.065 38.045 ;
        RECT 219.220 37.985 219.510 38.030 ;
        RECT 218.745 37.845 219.510 37.985 ;
        RECT 218.745 37.785 219.065 37.845 ;
        RECT 219.220 37.800 219.510 37.845 ;
        RECT 233.005 37.985 233.325 38.045 ;
        RECT 237.620 37.985 237.910 38.030 ;
        RECT 233.005 37.845 237.910 37.985 ;
        RECT 233.005 37.785 233.325 37.845 ;
        RECT 237.620 37.800 237.910 37.845 ;
        RECT 262.905 37.785 263.225 38.045 ;
        RECT 276.705 37.985 277.025 38.045 ;
        RECT 277.640 37.985 277.930 38.030 ;
        RECT 276.705 37.845 277.930 37.985 ;
        RECT 276.705 37.785 277.025 37.845 ;
        RECT 277.640 37.800 277.930 37.845 ;
        RECT 280.385 37.985 280.705 38.045 ;
        RECT 282.685 37.985 283.005 38.045 ;
        RECT 280.385 37.845 283.005 37.985 ;
        RECT 170.920 37.645 171.210 37.690 ;
        RECT 170.535 37.505 171.210 37.645 ;
        RECT 170.535 37.350 170.675 37.505 ;
        RECT 170.920 37.460 171.210 37.505 ;
        RECT 185.130 37.645 185.420 37.690 ;
        RECT 187.020 37.645 187.310 37.690 ;
        RECT 190.140 37.645 190.430 37.690 ;
        RECT 204.500 37.645 204.790 37.690 ;
        RECT 229.750 37.645 230.040 37.690 ;
        RECT 231.640 37.645 231.930 37.690 ;
        RECT 234.760 37.645 235.050 37.690 ;
        RECT 185.130 37.505 190.430 37.645 ;
        RECT 185.130 37.460 185.420 37.505 ;
        RECT 187.020 37.460 187.310 37.505 ;
        RECT 190.140 37.460 190.430 37.505 ;
        RECT 197.675 37.505 204.790 37.645 ;
        RECT 170.460 37.120 170.750 37.350 ;
        RECT 174.140 37.305 174.430 37.350 ;
        RECT 178.280 37.305 178.570 37.350 ;
        RECT 174.140 37.165 178.570 37.305 ;
        RECT 174.140 37.120 174.430 37.165 ;
        RECT 178.280 37.120 178.570 37.165 ;
        RECT 172.760 36.625 173.050 36.670 ;
        RECT 175.965 36.625 176.285 36.685 ;
        RECT 172.760 36.485 176.285 36.625 ;
        RECT 172.760 36.440 173.050 36.485 ;
        RECT 175.965 36.425 176.285 36.485 ;
        RECT 176.425 36.625 176.745 36.685 ;
        RECT 177.820 36.625 178.110 36.670 ;
        RECT 176.425 36.485 178.110 36.625 ;
        RECT 178.355 36.625 178.495 37.120 ;
        RECT 185.625 37.105 185.945 37.365 ;
        RECT 197.675 37.350 197.815 37.505 ;
        RECT 204.500 37.460 204.790 37.505 ;
        RECT 207.335 37.505 218.515 37.645 ;
        RECT 197.600 37.120 197.890 37.350 ;
        RECT 198.505 37.305 198.825 37.365 ;
        RECT 207.335 37.350 207.475 37.505 ;
        RECT 207.260 37.305 207.550 37.350 ;
        RECT 198.505 37.165 207.550 37.305 ;
        RECT 198.505 37.105 198.825 37.165 ;
        RECT 207.260 37.120 207.550 37.165 ;
        RECT 211.860 37.305 212.150 37.350 ;
        RECT 215.525 37.305 215.845 37.365 ;
        RECT 218.375 37.350 218.515 37.505 ;
        RECT 229.750 37.505 235.050 37.645 ;
        RECT 229.750 37.460 230.040 37.505 ;
        RECT 231.640 37.460 231.930 37.505 ;
        RECT 234.760 37.460 235.050 37.505 ;
        RECT 240.790 37.645 241.080 37.690 ;
        RECT 242.680 37.645 242.970 37.690 ;
        RECT 245.800 37.645 246.090 37.690 ;
        RECT 240.790 37.505 246.090 37.645 ;
        RECT 240.790 37.460 241.080 37.505 ;
        RECT 242.680 37.460 242.970 37.505 ;
        RECT 245.800 37.460 246.090 37.505 ;
        RECT 255.050 37.645 255.340 37.690 ;
        RECT 256.940 37.645 257.230 37.690 ;
        RECT 260.060 37.645 260.350 37.690 ;
        RECT 255.050 37.505 260.350 37.645 ;
        RECT 255.050 37.460 255.340 37.505 ;
        RECT 256.940 37.460 257.230 37.505 ;
        RECT 260.060 37.460 260.350 37.505 ;
        RECT 262.445 37.645 262.765 37.705 ;
        RECT 263.380 37.645 263.670 37.690 ;
        RECT 262.445 37.505 263.670 37.645 ;
        RECT 262.445 37.445 262.765 37.505 ;
        RECT 263.380 37.460 263.670 37.505 ;
        RECT 269.770 37.645 270.060 37.690 ;
        RECT 271.660 37.645 271.950 37.690 ;
        RECT 274.780 37.645 275.070 37.690 ;
        RECT 269.770 37.505 275.070 37.645 ;
        RECT 277.715 37.645 277.855 37.800 ;
        RECT 280.385 37.785 280.705 37.845 ;
        RECT 282.685 37.785 283.005 37.845 ;
        RECT 278.560 37.645 278.850 37.690 ;
        RECT 277.715 37.505 278.850 37.645 ;
        RECT 269.770 37.460 270.060 37.505 ;
        RECT 271.660 37.460 271.950 37.505 ;
        RECT 274.780 37.460 275.070 37.505 ;
        RECT 278.560 37.460 278.850 37.505 ;
        RECT 281.305 37.445 281.625 37.705 ;
        RECT 307.525 37.645 307.845 37.705 ;
        RECT 308.000 37.645 308.290 37.690 ;
        RECT 307.525 37.505 308.290 37.645 ;
        RECT 307.525 37.445 307.845 37.505 ;
        RECT 308.000 37.460 308.290 37.505 ;
        RECT 211.860 37.165 215.845 37.305 ;
        RECT 211.860 37.120 212.150 37.165 ;
        RECT 215.525 37.105 215.845 37.165 ;
        RECT 218.300 37.305 218.590 37.350 ;
        RECT 221.045 37.305 221.365 37.365 ;
        RECT 218.300 37.165 221.365 37.305 ;
        RECT 218.300 37.120 218.590 37.165 ;
        RECT 221.045 37.105 221.365 37.165 ;
        RECT 222.440 37.305 222.730 37.350 ;
        RECT 222.885 37.305 223.205 37.365 ;
        RECT 222.440 37.165 223.205 37.305 ;
        RECT 222.440 37.120 222.730 37.165 ;
        RECT 222.885 37.105 223.205 37.165 ;
        RECT 223.805 37.305 224.125 37.365 ;
        RECT 228.880 37.305 229.170 37.350 ;
        RECT 223.805 37.165 229.170 37.305 ;
        RECT 223.805 37.105 224.125 37.165 ;
        RECT 228.880 37.120 229.170 37.165 ;
        RECT 230.245 37.105 230.565 37.365 ;
        RECT 239.920 37.305 240.210 37.350 ;
        RECT 244.505 37.305 244.825 37.365 ;
        RECT 239.920 37.165 244.825 37.305 ;
        RECT 239.920 37.120 240.210 37.165 ;
        RECT 244.505 37.105 244.825 37.165 ;
        RECT 254.180 37.305 254.470 37.350 ;
        RECT 256.005 37.305 256.325 37.365 ;
        RECT 268.900 37.305 269.190 37.350 ;
        RECT 254.180 37.165 269.190 37.305 ;
        RECT 254.180 37.120 254.470 37.165 ;
        RECT 256.005 37.105 256.325 37.165 ;
        RECT 268.900 37.120 269.190 37.165 ;
        RECT 270.280 37.305 270.570 37.350 ;
        RECT 278.085 37.305 278.405 37.365 ;
        RECT 270.280 37.165 278.405 37.305 ;
        RECT 270.280 37.120 270.570 37.165 ;
        RECT 278.085 37.105 278.405 37.165 ;
        RECT 178.725 36.965 179.045 37.025 ;
        RECT 180.580 36.965 180.870 37.010 ;
        RECT 178.725 36.825 180.870 36.965 ;
        RECT 178.725 36.765 179.045 36.825 ;
        RECT 180.580 36.780 180.870 36.825 ;
        RECT 184.245 36.765 184.565 37.025 ;
        RECT 184.725 36.965 185.015 37.010 ;
        RECT 186.560 36.965 186.850 37.010 ;
        RECT 190.140 36.965 190.430 37.010 ;
        RECT 184.725 36.825 190.430 36.965 ;
        RECT 184.725 36.780 185.015 36.825 ;
        RECT 186.560 36.780 186.850 36.825 ;
        RECT 190.140 36.780 190.430 36.825 ;
        RECT 191.220 36.965 191.510 36.985 ;
        RECT 192.985 36.965 193.305 37.025 ;
        RECT 191.220 36.825 193.305 36.965 ;
        RECT 191.220 36.670 191.510 36.825 ;
        RECT 192.985 36.765 193.305 36.825 ;
        RECT 196.205 36.765 196.525 37.025 ;
        RECT 187.920 36.625 188.570 36.670 ;
        RECT 191.220 36.625 191.810 36.670 ;
        RECT 193.905 36.625 194.225 36.685 ;
        RECT 198.595 36.625 198.735 37.105 ;
        RECT 216.920 36.965 217.210 37.010 ;
        RECT 218.745 36.965 219.065 37.025 ;
        RECT 216.920 36.825 219.065 36.965 ;
        RECT 216.920 36.780 217.210 36.825 ;
        RECT 218.745 36.765 219.065 36.825 ;
        RECT 225.645 36.765 225.965 37.025 ;
        RECT 229.345 36.965 229.635 37.010 ;
        RECT 231.180 36.965 231.470 37.010 ;
        RECT 234.760 36.965 235.050 37.010 ;
        RECT 229.345 36.825 235.050 36.965 ;
        RECT 229.345 36.780 229.635 36.825 ;
        RECT 231.180 36.780 231.470 36.825 ;
        RECT 234.760 36.780 235.050 36.825 ;
        RECT 178.355 36.485 185.395 36.625 ;
        RECT 176.425 36.425 176.745 36.485 ;
        RECT 177.820 36.440 178.110 36.485 ;
        RECT 185.255 36.345 185.395 36.485 ;
        RECT 187.920 36.485 191.810 36.625 ;
        RECT 187.920 36.440 188.570 36.485 ;
        RECT 191.520 36.440 191.810 36.485 ;
        RECT 192.155 36.485 198.735 36.625 ;
        RECT 206.340 36.625 206.630 36.670 ;
        RECT 208.625 36.625 208.945 36.685 ;
        RECT 206.340 36.485 208.945 36.625 ;
        RECT 173.220 36.285 173.510 36.330 ;
        RECT 174.585 36.285 174.905 36.345 ;
        RECT 173.220 36.145 174.905 36.285 ;
        RECT 173.220 36.100 173.510 36.145 ;
        RECT 174.585 36.085 174.905 36.145 ;
        RECT 177.360 36.285 177.650 36.330 ;
        RECT 180.565 36.285 180.885 36.345 ;
        RECT 177.360 36.145 180.885 36.285 ;
        RECT 177.360 36.100 177.650 36.145 ;
        RECT 180.565 36.085 180.885 36.145 ;
        RECT 185.165 36.285 185.485 36.345 ;
        RECT 192.155 36.285 192.295 36.485 ;
        RECT 193.905 36.425 194.225 36.485 ;
        RECT 206.340 36.440 206.630 36.485 ;
        RECT 208.625 36.425 208.945 36.485 ;
        RECT 212.780 36.625 213.070 36.670 ;
        RECT 216.445 36.625 216.765 36.685 ;
        RECT 235.840 36.670 236.130 36.985 ;
        RECT 240.385 36.965 240.675 37.010 ;
        RECT 242.220 36.965 242.510 37.010 ;
        RECT 245.800 36.965 246.090 37.010 ;
        RECT 240.385 36.825 246.090 36.965 ;
        RECT 240.385 36.780 240.675 36.825 ;
        RECT 242.220 36.780 242.510 36.825 ;
        RECT 245.800 36.780 246.090 36.825 ;
        RECT 212.780 36.485 216.765 36.625 ;
        RECT 212.780 36.440 213.070 36.485 ;
        RECT 216.445 36.425 216.765 36.485 ;
        RECT 232.540 36.625 233.190 36.670 ;
        RECT 235.840 36.625 236.430 36.670 ;
        RECT 236.685 36.625 237.005 36.685 ;
        RECT 232.540 36.485 237.005 36.625 ;
        RECT 232.540 36.440 233.190 36.485 ;
        RECT 236.140 36.440 236.430 36.485 ;
        RECT 236.685 36.425 237.005 36.485 ;
        RECT 241.285 36.425 241.605 36.685 ;
        RECT 244.045 36.670 244.365 36.685 ;
        RECT 243.580 36.625 244.365 36.670 ;
        RECT 246.880 36.670 247.170 36.985 ;
        RECT 254.645 36.965 254.935 37.010 ;
        RECT 256.480 36.965 256.770 37.010 ;
        RECT 260.060 36.965 260.350 37.010 ;
        RECT 254.645 36.825 260.350 36.965 ;
        RECT 254.645 36.780 254.935 36.825 ;
        RECT 256.480 36.780 256.770 36.825 ;
        RECT 260.060 36.780 260.350 36.825 ;
        RECT 246.880 36.625 247.470 36.670 ;
        RECT 243.580 36.485 247.470 36.625 ;
        RECT 243.580 36.440 244.365 36.485 ;
        RECT 247.180 36.440 247.470 36.485 ;
        RECT 255.560 36.625 255.850 36.670 ;
        RECT 256.925 36.625 257.245 36.685 ;
        RECT 261.140 36.670 261.430 36.985 ;
        RECT 262.905 36.965 263.225 37.025 ;
        RECT 264.300 36.965 264.590 37.010 ;
        RECT 262.905 36.825 264.590 36.965 ;
        RECT 262.905 36.765 263.225 36.825 ;
        RECT 264.300 36.780 264.590 36.825 ;
        RECT 266.585 36.765 266.905 37.025 ;
        RECT 267.045 36.765 267.365 37.025 ;
        RECT 269.365 36.965 269.655 37.010 ;
        RECT 271.200 36.965 271.490 37.010 ;
        RECT 274.780 36.965 275.070 37.010 ;
        RECT 269.365 36.825 275.070 36.965 ;
        RECT 269.365 36.780 269.655 36.825 ;
        RECT 271.200 36.780 271.490 36.825 ;
        RECT 274.780 36.780 275.070 36.825 ;
        RECT 275.860 36.670 276.150 36.985 ;
        RECT 257.840 36.625 258.490 36.670 ;
        RECT 261.140 36.625 261.730 36.670 ;
        RECT 255.560 36.485 257.245 36.625 ;
        RECT 255.560 36.440 255.850 36.485 ;
        RECT 244.045 36.425 244.365 36.440 ;
        RECT 256.925 36.425 257.245 36.485 ;
        RECT 257.475 36.485 261.730 36.625 ;
        RECT 185.165 36.145 192.295 36.285 ;
        RECT 185.165 36.085 185.485 36.145 ;
        RECT 193.445 36.085 193.765 36.345 ;
        RECT 200.360 36.285 200.650 36.330 ;
        RECT 202.645 36.285 202.965 36.345 ;
        RECT 200.360 36.145 202.965 36.285 ;
        RECT 200.360 36.100 200.650 36.145 ;
        RECT 202.645 36.085 202.965 36.145 ;
        RECT 206.785 36.085 207.105 36.345 ;
        RECT 212.305 36.085 212.625 36.345 ;
        RECT 214.605 36.085 214.925 36.345 ;
        RECT 217.365 36.085 217.685 36.345 ;
        RECT 222.900 36.285 223.190 36.330 ;
        RECT 225.645 36.285 225.965 36.345 ;
        RECT 222.900 36.145 225.965 36.285 ;
        RECT 222.900 36.100 223.190 36.145 ;
        RECT 225.645 36.085 225.965 36.145 ;
        RECT 245.425 36.285 245.745 36.345 ;
        RECT 248.660 36.285 248.950 36.330 ;
        RECT 245.425 36.145 248.950 36.285 ;
        RECT 245.425 36.085 245.745 36.145 ;
        RECT 248.660 36.100 248.950 36.145 ;
        RECT 255.085 36.285 255.405 36.345 ;
        RECT 257.475 36.285 257.615 36.485 ;
        RECT 257.840 36.440 258.490 36.485 ;
        RECT 261.440 36.440 261.730 36.485 ;
        RECT 265.220 36.625 265.510 36.670 ;
        RECT 272.560 36.625 273.210 36.670 ;
        RECT 275.860 36.625 276.450 36.670 ;
        RECT 279.465 36.625 279.785 36.685 ;
        RECT 265.220 36.485 265.620 36.625 ;
        RECT 272.560 36.485 279.785 36.625 ;
        RECT 265.220 36.440 265.510 36.485 ;
        RECT 272.560 36.440 273.210 36.485 ;
        RECT 276.160 36.440 276.450 36.485 ;
        RECT 255.085 36.145 257.615 36.285 ;
        RECT 259.225 36.285 259.545 36.345 ;
        RECT 265.295 36.285 265.435 36.440 ;
        RECT 279.465 36.425 279.785 36.485 ;
        RECT 280.400 36.625 280.690 36.670 ;
        RECT 280.845 36.625 281.165 36.685 ;
        RECT 280.400 36.485 281.165 36.625 ;
        RECT 280.400 36.440 280.690 36.485 ;
        RECT 280.845 36.425 281.165 36.485 ;
        RECT 308.905 36.425 309.225 36.685 ;
        RECT 265.680 36.285 265.970 36.330 ;
        RECT 259.225 36.145 265.970 36.285 ;
        RECT 255.085 36.085 255.405 36.145 ;
        RECT 259.225 36.085 259.545 36.145 ;
        RECT 265.680 36.100 265.970 36.145 ;
        RECT 162.095 35.465 311.135 35.945 ;
        RECT 175.060 35.265 175.350 35.310 ;
        RECT 175.965 35.265 176.285 35.325 ;
        RECT 175.060 35.125 176.285 35.265 ;
        RECT 175.060 35.080 175.350 35.125 ;
        RECT 175.965 35.065 176.285 35.125 ;
        RECT 178.725 35.065 179.045 35.325 ;
        RECT 193.445 35.265 193.765 35.325 ;
        RECT 189.855 35.125 193.765 35.265 ;
        RECT 183.785 34.970 184.105 34.985 ;
        RECT 169.520 34.925 170.170 34.970 ;
        RECT 173.120 34.925 173.410 34.970 ;
        RECT 169.520 34.785 173.410 34.925 ;
        RECT 169.520 34.740 170.170 34.785 ;
        RECT 172.820 34.740 173.410 34.785 ;
        RECT 180.220 34.925 180.510 34.970 ;
        RECT 183.460 34.925 184.110 34.970 ;
        RECT 186.545 34.925 186.865 34.985 ;
        RECT 189.855 34.970 189.995 35.125 ;
        RECT 193.445 35.065 193.765 35.125 ;
        RECT 198.045 35.265 198.365 35.325 ;
        RECT 199.885 35.265 200.205 35.325 ;
        RECT 210.940 35.265 211.230 35.310 ;
        RECT 233.020 35.265 233.310 35.310 ;
        RECT 233.465 35.265 233.785 35.325 ;
        RECT 198.045 35.125 211.230 35.265 ;
        RECT 198.045 35.065 198.365 35.125 ;
        RECT 199.885 35.065 200.205 35.125 ;
        RECT 210.940 35.080 211.230 35.125 ;
        RECT 216.075 35.125 220.815 35.265 ;
        RECT 180.220 34.785 186.865 34.925 ;
        RECT 180.220 34.740 180.810 34.785 ;
        RECT 183.460 34.740 184.110 34.785 ;
        RECT 172.820 34.645 173.110 34.740 ;
        RECT 165.845 34.385 166.165 34.645 ;
        RECT 166.325 34.585 166.615 34.630 ;
        RECT 168.160 34.585 168.450 34.630 ;
        RECT 171.740 34.585 172.030 34.630 ;
        RECT 166.325 34.445 172.030 34.585 ;
        RECT 166.325 34.400 166.615 34.445 ;
        RECT 168.160 34.400 168.450 34.445 ;
        RECT 171.740 34.400 172.030 34.445 ;
        RECT 172.745 34.425 173.110 34.645 ;
        RECT 176.885 34.585 177.205 34.645 ;
        RECT 177.820 34.585 178.110 34.630 ;
        RECT 176.885 34.445 178.110 34.585 ;
        RECT 172.745 34.385 173.065 34.425 ;
        RECT 176.885 34.385 177.205 34.445 ;
        RECT 177.820 34.400 178.110 34.445 ;
        RECT 180.520 34.425 180.810 34.740 ;
        RECT 183.785 34.725 184.105 34.740 ;
        RECT 186.545 34.725 186.865 34.785 ;
        RECT 189.780 34.740 190.070 34.970 ;
        RECT 192.060 34.925 192.710 34.970 ;
        RECT 195.660 34.925 195.950 34.970 ;
        RECT 198.505 34.925 198.825 34.985 ;
        RECT 192.060 34.785 198.825 34.925 ;
        RECT 192.060 34.740 192.710 34.785 ;
        RECT 195.360 34.740 195.950 34.785 ;
        RECT 181.600 34.585 181.890 34.630 ;
        RECT 185.180 34.585 185.470 34.630 ;
        RECT 187.015 34.585 187.305 34.630 ;
        RECT 181.600 34.445 187.305 34.585 ;
        RECT 181.600 34.400 181.890 34.445 ;
        RECT 185.180 34.400 185.470 34.445 ;
        RECT 187.015 34.400 187.305 34.445 ;
        RECT 187.465 34.585 187.785 34.645 ;
        RECT 188.400 34.585 188.690 34.630 ;
        RECT 187.465 34.445 188.690 34.585 ;
        RECT 187.465 34.385 187.785 34.445 ;
        RECT 188.400 34.400 188.690 34.445 ;
        RECT 188.865 34.585 189.155 34.630 ;
        RECT 190.700 34.585 190.990 34.630 ;
        RECT 194.280 34.585 194.570 34.630 ;
        RECT 188.865 34.445 194.570 34.585 ;
        RECT 188.865 34.400 189.155 34.445 ;
        RECT 190.700 34.400 190.990 34.445 ;
        RECT 194.280 34.400 194.570 34.445 ;
        RECT 195.360 34.425 195.650 34.740 ;
        RECT 198.505 34.725 198.825 34.785 ;
        RECT 202.645 34.725 202.965 34.985 ;
        RECT 204.940 34.925 205.590 34.970 ;
        RECT 208.540 34.925 208.830 34.970 ;
        RECT 209.085 34.925 209.405 34.985 ;
        RECT 216.075 34.925 216.215 35.125 ;
        RECT 204.940 34.785 216.215 34.925 ;
        RECT 216.560 34.925 216.850 34.970 ;
        RECT 219.800 34.925 220.450 34.970 ;
        RECT 220.675 34.925 220.815 35.125 ;
        RECT 233.020 35.125 233.785 35.265 ;
        RECT 233.020 35.080 233.310 35.125 ;
        RECT 233.465 35.065 233.785 35.125 ;
        RECT 236.240 35.265 236.530 35.310 ;
        RECT 236.685 35.265 237.005 35.325 ;
        RECT 249.120 35.265 249.410 35.310 ;
        RECT 252.325 35.265 252.645 35.325 ;
        RECT 255.085 35.265 255.405 35.325 ;
        RECT 262.920 35.265 263.210 35.310 ;
        RECT 267.045 35.265 267.365 35.325 ;
        RECT 236.240 35.125 237.005 35.265 ;
        RECT 236.240 35.080 236.530 35.125 ;
        RECT 221.965 34.925 222.285 34.985 ;
        RECT 216.560 34.785 222.285 34.925 ;
        RECT 204.940 34.740 205.590 34.785 ;
        RECT 208.240 34.740 208.830 34.785 ;
        RECT 200.805 34.585 201.125 34.645 ;
        RECT 201.280 34.585 201.570 34.630 ;
        RECT 200.805 34.445 201.570 34.585 ;
        RECT 200.805 34.385 201.125 34.445 ;
        RECT 201.280 34.400 201.570 34.445 ;
        RECT 201.745 34.585 202.035 34.630 ;
        RECT 203.580 34.585 203.870 34.630 ;
        RECT 207.160 34.585 207.450 34.630 ;
        RECT 201.745 34.445 207.450 34.585 ;
        RECT 201.745 34.400 202.035 34.445 ;
        RECT 203.580 34.400 203.870 34.445 ;
        RECT 207.160 34.400 207.450 34.445 ;
        RECT 208.240 34.425 208.530 34.740 ;
        RECT 209.085 34.725 209.405 34.785 ;
        RECT 216.560 34.740 217.150 34.785 ;
        RECT 219.800 34.740 220.450 34.785 ;
        RECT 212.320 34.585 212.610 34.630 ;
        RECT 212.765 34.585 213.085 34.645 ;
        RECT 212.320 34.445 213.085 34.585 ;
        RECT 212.320 34.400 212.610 34.445 ;
        RECT 212.765 34.385 213.085 34.445 ;
        RECT 216.860 34.425 217.150 34.740 ;
        RECT 221.965 34.725 222.285 34.785 ;
        RECT 225.645 34.725 225.965 34.985 ;
        RECT 227.940 34.925 228.590 34.970 ;
        RECT 231.540 34.925 231.830 34.970 ;
        RECT 236.315 34.925 236.455 35.080 ;
        RECT 236.685 35.065 237.005 35.125 ;
        RECT 243.675 35.125 248.875 35.265 ;
        RECT 227.940 34.785 236.455 34.925 ;
        RECT 241.760 34.925 242.050 34.970 ;
        RECT 242.205 34.925 242.525 34.985 ;
        RECT 241.760 34.785 242.525 34.925 ;
        RECT 243.675 34.925 243.815 35.125 ;
        RECT 244.045 34.970 244.365 34.985 ;
        RECT 244.040 34.925 244.690 34.970 ;
        RECT 247.640 34.925 247.930 34.970 ;
        RECT 243.675 34.785 247.930 34.925 ;
        RECT 248.735 34.925 248.875 35.125 ;
        RECT 249.120 35.125 252.645 35.265 ;
        RECT 249.120 35.080 249.410 35.125 ;
        RECT 252.325 35.065 252.645 35.125 ;
        RECT 253.795 35.125 256.695 35.265 ;
        RECT 253.795 34.925 253.935 35.125 ;
        RECT 255.085 35.065 255.405 35.125 ;
        RECT 256.005 34.925 256.325 34.985 ;
        RECT 248.735 34.785 253.935 34.925 ;
        RECT 254.255 34.785 256.325 34.925 ;
        RECT 256.555 34.925 256.695 35.125 ;
        RECT 262.920 35.125 267.365 35.265 ;
        RECT 262.920 35.080 263.210 35.125 ;
        RECT 267.045 35.065 267.365 35.125 ;
        RECT 280.385 35.065 280.705 35.325 ;
        RECT 257.840 34.925 258.490 34.970 ;
        RECT 261.440 34.925 261.730 34.970 ;
        RECT 256.555 34.785 261.730 34.925 ;
        RECT 227.940 34.740 228.590 34.785 ;
        RECT 231.240 34.740 231.830 34.785 ;
        RECT 241.760 34.740 242.050 34.785 ;
        RECT 217.940 34.585 218.230 34.630 ;
        RECT 221.520 34.585 221.810 34.630 ;
        RECT 223.355 34.585 223.645 34.630 ;
        RECT 217.940 34.445 223.645 34.585 ;
        RECT 217.940 34.400 218.230 34.445 ;
        RECT 221.520 34.400 221.810 34.445 ;
        RECT 223.355 34.400 223.645 34.445 ;
        RECT 224.745 34.585 225.035 34.630 ;
        RECT 226.580 34.585 226.870 34.630 ;
        RECT 230.160 34.585 230.450 34.630 ;
        RECT 224.745 34.445 230.450 34.585 ;
        RECT 224.745 34.400 225.035 34.445 ;
        RECT 226.580 34.400 226.870 34.445 ;
        RECT 230.160 34.400 230.450 34.445 ;
        RECT 231.240 34.425 231.530 34.740 ;
        RECT 242.205 34.725 242.525 34.785 ;
        RECT 244.040 34.740 244.690 34.785 ;
        RECT 247.340 34.740 247.930 34.785 ;
        RECT 244.045 34.725 244.365 34.740 ;
        RECT 232.545 34.585 232.865 34.645 ;
        RECT 236.700 34.585 236.990 34.630 ;
        RECT 232.545 34.445 236.990 34.585 ;
        RECT 232.545 34.385 232.865 34.445 ;
        RECT 236.700 34.400 236.990 34.445 ;
        RECT 240.845 34.585 241.135 34.630 ;
        RECT 242.680 34.585 242.970 34.630 ;
        RECT 246.260 34.585 246.550 34.630 ;
        RECT 240.845 34.445 246.550 34.585 ;
        RECT 240.845 34.400 241.135 34.445 ;
        RECT 242.680 34.400 242.970 34.445 ;
        RECT 246.260 34.400 246.550 34.445 ;
        RECT 247.340 34.425 247.630 34.740 ;
        RECT 248.185 34.585 248.505 34.645 ;
        RECT 254.255 34.630 254.395 34.785 ;
        RECT 256.005 34.725 256.325 34.785 ;
        RECT 257.840 34.740 258.490 34.785 ;
        RECT 261.140 34.740 261.730 34.785 ;
        RECT 254.180 34.585 254.470 34.630 ;
        RECT 248.185 34.445 254.470 34.585 ;
        RECT 248.185 34.385 248.505 34.445 ;
        RECT 254.180 34.400 254.470 34.445 ;
        RECT 254.645 34.585 254.935 34.630 ;
        RECT 256.480 34.585 256.770 34.630 ;
        RECT 260.060 34.585 260.350 34.630 ;
        RECT 254.645 34.445 260.350 34.585 ;
        RECT 254.645 34.400 254.935 34.445 ;
        RECT 256.480 34.400 256.770 34.445 ;
        RECT 260.060 34.400 260.350 34.445 ;
        RECT 261.140 34.425 261.430 34.740 ;
        RECT 273.025 34.725 273.345 34.985 ;
        RECT 275.320 34.925 275.970 34.970 ;
        RECT 278.920 34.925 279.210 34.970 ;
        RECT 279.465 34.925 279.785 34.985 ;
        RECT 283.145 34.925 283.465 34.985 ;
        RECT 275.320 34.785 283.465 34.925 ;
        RECT 275.320 34.740 275.970 34.785 ;
        RECT 278.620 34.740 279.210 34.785 ;
        RECT 271.645 34.385 271.965 34.645 ;
        RECT 272.125 34.585 272.415 34.630 ;
        RECT 273.960 34.585 274.250 34.630 ;
        RECT 277.540 34.585 277.830 34.630 ;
        RECT 272.125 34.445 277.830 34.585 ;
        RECT 272.125 34.400 272.415 34.445 ;
        RECT 273.960 34.400 274.250 34.445 ;
        RECT 277.540 34.400 277.830 34.445 ;
        RECT 278.620 34.425 278.910 34.740 ;
        RECT 279.465 34.725 279.785 34.785 ;
        RECT 283.145 34.725 283.465 34.785 ;
        RECT 167.240 34.245 167.530 34.290 ;
        RECT 170.905 34.245 171.225 34.305 ;
        RECT 167.240 34.105 171.225 34.245 ;
        RECT 167.240 34.060 167.530 34.105 ;
        RECT 170.905 34.045 171.225 34.105 ;
        RECT 186.085 34.045 186.405 34.305 ;
        RECT 197.140 34.245 197.430 34.290 ;
        RECT 200.360 34.245 200.650 34.290 ;
        RECT 197.140 34.105 200.650 34.245 ;
        RECT 197.140 34.060 197.430 34.105 ;
        RECT 200.360 34.060 200.650 34.105 ;
        RECT 222.425 34.045 222.745 34.305 ;
        RECT 223.805 34.245 224.125 34.305 ;
        RECT 224.280 34.245 224.570 34.290 ;
        RECT 223.805 34.105 224.570 34.245 ;
        RECT 223.805 34.045 224.125 34.105 ;
        RECT 224.280 34.060 224.570 34.105 ;
        RECT 240.380 34.060 240.670 34.290 ;
        RECT 242.205 34.245 242.525 34.305 ;
        RECT 244.965 34.245 245.285 34.305 ;
        RECT 242.205 34.105 245.285 34.245 ;
        RECT 166.730 33.905 167.020 33.950 ;
        RECT 168.620 33.905 168.910 33.950 ;
        RECT 171.740 33.905 172.030 33.950 ;
        RECT 166.730 33.765 172.030 33.905 ;
        RECT 166.730 33.720 167.020 33.765 ;
        RECT 168.620 33.720 168.910 33.765 ;
        RECT 171.740 33.720 172.030 33.765 ;
        RECT 174.600 33.905 174.890 33.950 ;
        RECT 175.965 33.905 176.285 33.965 ;
        RECT 174.600 33.765 176.285 33.905 ;
        RECT 174.600 33.720 174.890 33.765 ;
        RECT 175.965 33.705 176.285 33.765 ;
        RECT 181.600 33.905 181.890 33.950 ;
        RECT 184.720 33.905 185.010 33.950 ;
        RECT 186.610 33.905 186.900 33.950 ;
        RECT 181.600 33.765 186.900 33.905 ;
        RECT 181.600 33.720 181.890 33.765 ;
        RECT 184.720 33.720 185.010 33.765 ;
        RECT 186.610 33.720 186.900 33.765 ;
        RECT 189.270 33.905 189.560 33.950 ;
        RECT 191.160 33.905 191.450 33.950 ;
        RECT 194.280 33.905 194.570 33.950 ;
        RECT 189.270 33.765 194.570 33.905 ;
        RECT 189.270 33.720 189.560 33.765 ;
        RECT 191.160 33.720 191.450 33.765 ;
        RECT 194.280 33.720 194.570 33.765 ;
        RECT 202.150 33.905 202.440 33.950 ;
        RECT 204.040 33.905 204.330 33.950 ;
        RECT 207.160 33.905 207.450 33.950 ;
        RECT 202.150 33.765 207.450 33.905 ;
        RECT 202.150 33.720 202.440 33.765 ;
        RECT 204.040 33.720 204.330 33.765 ;
        RECT 207.160 33.720 207.450 33.765 ;
        RECT 217.940 33.905 218.230 33.950 ;
        RECT 221.060 33.905 221.350 33.950 ;
        RECT 222.950 33.905 223.240 33.950 ;
        RECT 217.940 33.765 223.240 33.905 ;
        RECT 217.940 33.720 218.230 33.765 ;
        RECT 221.060 33.720 221.350 33.765 ;
        RECT 222.950 33.720 223.240 33.765 ;
        RECT 225.150 33.905 225.440 33.950 ;
        RECT 227.040 33.905 227.330 33.950 ;
        RECT 230.160 33.905 230.450 33.950 ;
        RECT 225.150 33.765 230.450 33.905 ;
        RECT 225.150 33.720 225.440 33.765 ;
        RECT 227.040 33.720 227.330 33.765 ;
        RECT 230.160 33.720 230.450 33.765 ;
        RECT 192.065 33.565 192.385 33.625 ;
        RECT 197.600 33.565 197.890 33.610 ;
        RECT 192.065 33.425 197.890 33.565 ;
        RECT 192.065 33.365 192.385 33.425 ;
        RECT 197.600 33.380 197.890 33.425 ;
        RECT 210.005 33.365 210.325 33.625 ;
        RECT 215.080 33.565 215.370 33.610 ;
        RECT 217.365 33.565 217.685 33.625 ;
        RECT 219.205 33.565 219.525 33.625 ;
        RECT 215.080 33.425 219.525 33.565 ;
        RECT 240.455 33.565 240.595 34.060 ;
        RECT 242.205 34.045 242.525 34.105 ;
        RECT 244.965 34.045 245.285 34.105 ;
        RECT 255.560 34.245 255.850 34.290 ;
        RECT 257.385 34.245 257.705 34.305 ;
        RECT 255.560 34.105 257.705 34.245 ;
        RECT 255.560 34.060 255.850 34.105 ;
        RECT 257.385 34.045 257.705 34.105 ;
        RECT 241.250 33.905 241.540 33.950 ;
        RECT 243.140 33.905 243.430 33.950 ;
        RECT 246.260 33.905 246.550 33.950 ;
        RECT 241.250 33.765 246.550 33.905 ;
        RECT 241.250 33.720 241.540 33.765 ;
        RECT 243.140 33.720 243.430 33.765 ;
        RECT 246.260 33.720 246.550 33.765 ;
        RECT 255.050 33.905 255.340 33.950 ;
        RECT 256.940 33.905 257.230 33.950 ;
        RECT 260.060 33.905 260.350 33.950 ;
        RECT 255.050 33.765 260.350 33.905 ;
        RECT 255.050 33.720 255.340 33.765 ;
        RECT 256.940 33.720 257.230 33.765 ;
        RECT 260.060 33.720 260.350 33.765 ;
        RECT 272.530 33.905 272.820 33.950 ;
        RECT 274.420 33.905 274.710 33.950 ;
        RECT 277.540 33.905 277.830 33.950 ;
        RECT 272.530 33.765 277.830 33.905 ;
        RECT 272.530 33.720 272.820 33.765 ;
        RECT 274.420 33.720 274.710 33.765 ;
        RECT 277.540 33.720 277.830 33.765 ;
        RECT 244.505 33.565 244.825 33.625 ;
        RECT 240.455 33.425 244.825 33.565 ;
        RECT 215.080 33.380 215.370 33.425 ;
        RECT 217.365 33.365 217.685 33.425 ;
        RECT 219.205 33.365 219.525 33.425 ;
        RECT 244.505 33.365 244.825 33.425 ;
        RECT 162.095 32.745 311.135 33.225 ;
        RECT 195.300 32.545 195.590 32.590 ;
        RECT 196.205 32.545 196.525 32.605 ;
        RECT 183.875 32.405 191.835 32.545 ;
        RECT 166.730 32.205 167.020 32.250 ;
        RECT 168.620 32.205 168.910 32.250 ;
        RECT 171.740 32.205 172.030 32.250 ;
        RECT 166.730 32.065 172.030 32.205 ;
        RECT 166.730 32.020 167.020 32.065 ;
        RECT 168.620 32.020 168.910 32.065 ;
        RECT 171.740 32.020 172.030 32.065 ;
        RECT 165.860 31.865 166.150 31.910 ;
        RECT 167.685 31.865 168.005 31.925 ;
        RECT 165.860 31.725 168.005 31.865 ;
        RECT 165.860 31.680 166.150 31.725 ;
        RECT 167.685 31.665 168.005 31.725 ;
        RECT 174.585 31.665 174.905 31.925 ;
        RECT 176.425 31.865 176.745 31.925 ;
        RECT 177.820 31.865 178.110 31.910 ;
        RECT 176.425 31.725 178.110 31.865 ;
        RECT 176.425 31.665 176.745 31.725 ;
        RECT 177.820 31.680 178.110 31.725 ;
        RECT 178.725 31.865 179.045 31.925 ;
        RECT 183.875 31.865 184.015 32.405 ;
        RECT 191.695 32.265 191.835 32.405 ;
        RECT 195.300 32.405 196.525 32.545 ;
        RECT 195.300 32.360 195.590 32.405 ;
        RECT 196.205 32.345 196.525 32.405 ;
        RECT 206.785 32.545 207.105 32.605 ;
        RECT 207.260 32.545 207.550 32.590 ;
        RECT 215.525 32.545 215.845 32.605 ;
        RECT 222.425 32.545 222.745 32.605 ;
        RECT 227.040 32.545 227.330 32.590 ;
        RECT 242.205 32.545 242.525 32.605 ;
        RECT 206.785 32.405 207.550 32.545 ;
        RECT 206.785 32.345 207.105 32.405 ;
        RECT 207.260 32.360 207.550 32.405 ;
        RECT 207.795 32.405 221.505 32.545 ;
        RECT 184.245 32.005 184.565 32.265 ;
        RECT 185.280 32.205 185.570 32.250 ;
        RECT 188.400 32.205 188.690 32.250 ;
        RECT 190.290 32.205 190.580 32.250 ;
        RECT 185.280 32.065 190.580 32.205 ;
        RECT 185.280 32.020 185.570 32.065 ;
        RECT 188.400 32.020 188.690 32.065 ;
        RECT 190.290 32.020 190.580 32.065 ;
        RECT 191.605 32.205 191.925 32.265 ;
        RECT 207.795 32.205 207.935 32.405 ;
        RECT 215.525 32.345 215.845 32.405 ;
        RECT 191.605 32.065 207.935 32.205 ;
        RECT 210.120 32.205 210.410 32.250 ;
        RECT 213.240 32.205 213.530 32.250 ;
        RECT 215.130 32.205 215.420 32.250 ;
        RECT 210.120 32.065 215.420 32.205 ;
        RECT 221.365 32.205 221.505 32.405 ;
        RECT 222.425 32.405 227.330 32.545 ;
        RECT 222.425 32.345 222.745 32.405 ;
        RECT 227.040 32.360 227.330 32.405 ;
        RECT 230.795 32.405 242.525 32.545 ;
        RECT 230.795 32.205 230.935 32.405 ;
        RECT 242.205 32.345 242.525 32.405 ;
        RECT 242.665 32.545 242.985 32.605 ;
        RECT 243.200 32.545 243.490 32.590 ;
        RECT 242.665 32.405 243.490 32.545 ;
        RECT 242.665 32.345 242.985 32.405 ;
        RECT 243.200 32.360 243.490 32.405 ;
        RECT 221.365 32.065 230.935 32.205 ;
        RECT 238.640 32.205 238.930 32.250 ;
        RECT 241.760 32.205 242.050 32.250 ;
        RECT 243.650 32.205 243.940 32.250 ;
        RECT 238.640 32.065 243.940 32.205 ;
        RECT 191.605 32.005 191.925 32.065 ;
        RECT 178.725 31.725 184.015 31.865 ;
        RECT 184.335 31.865 184.475 32.005 ;
        RECT 184.335 31.725 191.375 31.865 ;
        RECT 178.725 31.665 179.045 31.725 ;
        RECT 166.325 31.525 166.615 31.570 ;
        RECT 168.160 31.525 168.450 31.570 ;
        RECT 171.740 31.525 172.030 31.570 ;
        RECT 166.325 31.385 172.030 31.525 ;
        RECT 166.325 31.340 166.615 31.385 ;
        RECT 168.160 31.340 168.450 31.385 ;
        RECT 171.740 31.340 172.030 31.385 ;
        RECT 172.745 31.545 173.065 31.585 ;
        RECT 172.745 31.325 173.110 31.545 ;
        RECT 174.675 31.525 174.815 31.665 ;
        RECT 176.885 31.525 177.205 31.585 ;
        RECT 191.235 31.570 191.375 31.725 ;
        RECT 192.540 31.680 192.830 31.910 ;
        RECT 193.000 31.865 193.290 31.910 ;
        RECT 196.665 31.865 196.985 31.925 ;
        RECT 204.575 31.910 204.715 32.065 ;
        RECT 210.120 32.020 210.410 32.065 ;
        RECT 213.240 32.020 213.530 32.065 ;
        RECT 215.130 32.020 215.420 32.065 ;
        RECT 203.580 31.865 203.870 31.910 ;
        RECT 193.000 31.725 203.870 31.865 ;
        RECT 193.000 31.680 193.290 31.725 ;
        RECT 177.360 31.525 177.650 31.570 ;
        RECT 174.675 31.385 177.650 31.525 ;
        RECT 176.885 31.325 177.205 31.385 ;
        RECT 177.360 31.340 177.650 31.385 ;
        RECT 167.225 30.985 167.545 31.245 ;
        RECT 172.820 31.230 173.110 31.325 ;
        RECT 184.200 31.230 184.490 31.545 ;
        RECT 185.280 31.525 185.570 31.570 ;
        RECT 188.860 31.525 189.150 31.570 ;
        RECT 190.695 31.525 190.985 31.570 ;
        RECT 185.280 31.385 190.985 31.525 ;
        RECT 185.280 31.340 185.570 31.385 ;
        RECT 188.860 31.340 189.150 31.385 ;
        RECT 190.695 31.340 190.985 31.385 ;
        RECT 191.160 31.340 191.450 31.570 ;
        RECT 192.615 31.525 192.755 31.680 ;
        RECT 196.665 31.665 196.985 31.725 ;
        RECT 203.580 31.680 203.870 31.725 ;
        RECT 204.500 31.680 204.790 31.910 ;
        RECT 212.305 31.865 212.625 31.925 ;
        RECT 207.335 31.725 212.625 31.865 ;
        RECT 193.905 31.525 194.225 31.585 ;
        RECT 192.615 31.385 194.225 31.525 ;
        RECT 169.520 31.185 170.170 31.230 ;
        RECT 172.820 31.185 173.410 31.230 ;
        RECT 169.520 31.045 173.410 31.185 ;
        RECT 169.520 31.000 170.170 31.045 ;
        RECT 173.120 31.000 173.410 31.045 ;
        RECT 183.900 31.185 184.490 31.230 ;
        RECT 186.545 31.185 186.865 31.245 ;
        RECT 187.140 31.185 187.790 31.230 ;
        RECT 183.900 31.045 187.790 31.185 ;
        RECT 183.900 31.000 184.190 31.045 ;
        RECT 186.545 30.985 186.865 31.045 ;
        RECT 187.140 31.000 187.790 31.045 ;
        RECT 189.765 30.985 190.085 31.245 ;
        RECT 191.235 31.185 191.375 31.340 ;
        RECT 193.905 31.325 194.225 31.385 ;
        RECT 197.600 31.525 197.890 31.570 ;
        RECT 203.120 31.525 203.410 31.570 ;
        RECT 207.335 31.525 207.475 31.725 ;
        RECT 212.305 31.665 212.625 31.725 ;
        RECT 214.605 31.665 214.925 31.925 ;
        RECT 216.000 31.865 216.290 31.910 ;
        RECT 223.805 31.865 224.125 31.925 ;
        RECT 230.335 31.910 230.475 32.065 ;
        RECT 238.640 32.020 238.930 32.065 ;
        RECT 241.760 32.020 242.050 32.065 ;
        RECT 243.650 32.020 243.940 32.065 ;
        RECT 216.000 31.725 224.125 31.865 ;
        RECT 216.000 31.680 216.290 31.725 ;
        RECT 223.805 31.665 224.125 31.725 ;
        RECT 230.260 31.680 230.550 31.910 ;
        RECT 235.780 31.865 236.070 31.910 ;
        RECT 232.175 31.725 236.070 31.865 ;
        RECT 209.085 31.545 209.405 31.585 ;
        RECT 197.600 31.385 201.495 31.525 ;
        RECT 197.600 31.340 197.890 31.385 ;
        RECT 200.805 31.185 201.125 31.245 ;
        RECT 191.235 31.045 201.125 31.185 ;
        RECT 200.805 30.985 201.125 31.045 ;
        RECT 175.505 30.645 175.825 30.905 ;
        RECT 180.565 30.845 180.885 30.905 ;
        RECT 182.420 30.845 182.710 30.890 ;
        RECT 180.565 30.705 182.710 30.845 ;
        RECT 180.565 30.645 180.885 30.705 ;
        RECT 182.420 30.660 182.710 30.705 ;
        RECT 192.065 30.845 192.385 30.905 ;
        RECT 193.460 30.845 193.750 30.890 ;
        RECT 192.065 30.705 193.750 30.845 ;
        RECT 192.065 30.645 192.385 30.705 ;
        RECT 193.460 30.660 193.750 30.705 ;
        RECT 200.345 30.645 200.665 30.905 ;
        RECT 201.355 30.890 201.495 31.385 ;
        RECT 203.120 31.385 207.475 31.525 ;
        RECT 203.120 31.340 203.410 31.385 ;
        RECT 209.040 31.325 209.405 31.545 ;
        RECT 210.120 31.525 210.410 31.570 ;
        RECT 213.700 31.525 213.990 31.570 ;
        RECT 215.535 31.525 215.825 31.570 ;
        RECT 210.120 31.385 215.825 31.525 ;
        RECT 210.120 31.340 210.410 31.385 ;
        RECT 213.700 31.340 213.990 31.385 ;
        RECT 215.535 31.340 215.825 31.385 ;
        RECT 216.445 31.325 216.765 31.585 ;
        RECT 219.205 31.325 219.525 31.585 ;
        RECT 227.945 31.525 228.265 31.585 ;
        RECT 232.175 31.570 232.315 31.725 ;
        RECT 235.780 31.680 236.070 31.725 ;
        RECT 244.505 31.865 244.825 31.925 ;
        RECT 248.185 31.865 248.505 31.925 ;
        RECT 244.505 31.725 248.505 31.865 ;
        RECT 244.505 31.665 244.825 31.725 ;
        RECT 248.185 31.665 248.505 31.725 ;
        RECT 259.240 31.865 259.530 31.910 ;
        RECT 261.985 31.865 262.305 31.925 ;
        RECT 259.240 31.725 262.305 31.865 ;
        RECT 259.240 31.680 259.530 31.725 ;
        RECT 261.985 31.665 262.305 31.725 ;
        RECT 232.100 31.525 232.390 31.570 ;
        RECT 227.945 31.385 232.390 31.525 ;
        RECT 227.945 31.325 228.265 31.385 ;
        RECT 232.100 31.340 232.390 31.385 ;
        RECT 209.040 31.230 209.330 31.325 ;
        RECT 208.740 31.185 209.330 31.230 ;
        RECT 211.980 31.185 212.630 31.230 ;
        RECT 208.740 31.045 212.630 31.185 ;
        RECT 216.535 31.185 216.675 31.325 ;
        RECT 237.560 31.230 237.850 31.545 ;
        RECT 238.640 31.525 238.930 31.570 ;
        RECT 242.220 31.525 242.510 31.570 ;
        RECT 244.055 31.525 244.345 31.570 ;
        RECT 238.640 31.385 244.345 31.525 ;
        RECT 238.640 31.340 238.930 31.385 ;
        RECT 242.220 31.340 242.510 31.385 ;
        RECT 244.055 31.340 244.345 31.385 ;
        RECT 258.765 31.325 259.085 31.585 ;
        RECT 259.685 31.325 260.005 31.585 ;
        RECT 229.340 31.185 229.630 31.230 ;
        RECT 216.535 31.045 229.630 31.185 ;
        RECT 208.740 31.000 209.030 31.045 ;
        RECT 211.980 31.000 212.630 31.045 ;
        RECT 229.340 31.000 229.630 31.045 ;
        RECT 237.260 31.185 237.850 31.230 ;
        RECT 240.500 31.185 241.150 31.230 ;
        RECT 243.585 31.185 243.905 31.245 ;
        RECT 237.260 31.045 243.905 31.185 ;
        RECT 237.260 31.000 237.550 31.045 ;
        RECT 240.500 31.000 241.150 31.045 ;
        RECT 243.585 30.985 243.905 31.045 ;
        RECT 201.280 30.660 201.570 30.890 ;
        RECT 228.880 30.845 229.170 30.890 ;
        RECT 235.320 30.845 235.610 30.890 ;
        RECT 243.125 30.845 243.445 30.905 ;
        RECT 228.880 30.705 243.445 30.845 ;
        RECT 228.880 30.660 229.170 30.705 ;
        RECT 235.320 30.660 235.610 30.705 ;
        RECT 243.125 30.645 243.445 30.705 ;
        RECT 162.095 30.025 311.135 30.505 ;
        RECT 167.225 29.825 167.545 29.885 ;
        RECT 168.620 29.825 168.910 29.870 ;
        RECT 167.225 29.685 168.910 29.825 ;
        RECT 167.225 29.625 167.545 29.685 ;
        RECT 168.620 29.640 168.910 29.685 ;
        RECT 176.425 29.825 176.745 29.885 ;
        RECT 179.660 29.825 179.950 29.870 ;
        RECT 176.425 29.685 179.950 29.825 ;
        RECT 176.425 29.625 176.745 29.685 ;
        RECT 179.660 29.640 179.950 29.685 ;
        RECT 183.340 29.825 183.630 29.870 ;
        RECT 186.085 29.825 186.405 29.885 ;
        RECT 183.340 29.685 186.405 29.825 ;
        RECT 183.340 29.640 183.630 29.685 ;
        RECT 186.085 29.625 186.405 29.685 ;
        RECT 196.665 29.625 196.985 29.885 ;
        RECT 200.805 29.825 201.125 29.885 ;
        RECT 200.805 29.685 205.175 29.825 ;
        RECT 200.805 29.625 201.125 29.685 ;
        RECT 174.140 29.485 174.430 29.530 ;
        RECT 180.565 29.485 180.885 29.545 ;
        RECT 174.140 29.345 180.885 29.485 ;
        RECT 174.140 29.300 174.430 29.345 ;
        RECT 180.565 29.285 180.885 29.345 ;
        RECT 185.625 29.285 185.945 29.545 ;
        RECT 190.700 29.485 190.990 29.530 ;
        RECT 186.175 29.345 190.990 29.485 ;
        RECT 164.940 29.145 165.230 29.190 ;
        RECT 172.285 29.145 172.605 29.205 ;
        RECT 164.940 29.005 172.605 29.145 ;
        RECT 164.940 28.960 165.230 29.005 ;
        RECT 172.285 28.945 172.605 29.005 ;
        RECT 175.965 29.145 176.285 29.205 ;
        RECT 176.440 29.145 176.730 29.190 ;
        RECT 175.965 29.005 176.730 29.145 ;
        RECT 180.655 29.145 180.795 29.285 ;
        RECT 186.175 29.190 186.315 29.345 ;
        RECT 190.700 29.300 190.990 29.345 ;
        RECT 186.100 29.145 186.390 29.190 ;
        RECT 180.655 29.005 186.390 29.145 ;
        RECT 175.965 28.945 176.285 29.005 ;
        RECT 176.440 28.960 176.730 29.005 ;
        RECT 186.100 28.960 186.390 29.005 ;
        RECT 190.240 29.145 190.530 29.190 ;
        RECT 193.000 29.145 193.290 29.190 ;
        RECT 190.240 29.005 193.290 29.145 ;
        RECT 190.240 28.960 190.530 29.005 ;
        RECT 193.000 28.960 193.290 29.005 ;
        RECT 196.220 29.145 196.510 29.190 ;
        RECT 196.755 29.145 196.895 29.625 ;
        RECT 198.160 29.485 198.450 29.530 ;
        RECT 201.400 29.485 202.050 29.530 ;
        RECT 198.160 29.345 202.050 29.485 ;
        RECT 205.035 29.485 205.175 29.685 ;
        RECT 208.625 29.625 208.945 29.885 ;
        RECT 205.035 29.345 205.635 29.485 ;
        RECT 198.160 29.300 198.750 29.345 ;
        RECT 201.400 29.300 202.050 29.345 ;
        RECT 196.220 29.005 196.895 29.145 ;
        RECT 198.460 29.205 198.750 29.300 ;
        RECT 196.220 28.960 196.510 29.005 ;
        RECT 198.460 28.985 198.825 29.205 ;
        RECT 205.495 29.190 205.635 29.345 ;
        RECT 198.505 28.945 198.825 28.985 ;
        RECT 199.540 29.145 199.830 29.190 ;
        RECT 203.120 29.145 203.410 29.190 ;
        RECT 204.955 29.145 205.245 29.190 ;
        RECT 199.540 29.005 205.245 29.145 ;
        RECT 199.540 28.960 199.830 29.005 ;
        RECT 203.120 28.960 203.410 29.005 ;
        RECT 204.955 28.960 205.245 29.005 ;
        RECT 205.420 28.960 205.710 29.190 ;
        RECT 210.005 29.145 210.325 29.205 ;
        RECT 211.400 29.145 211.690 29.190 ;
        RECT 210.005 29.005 211.690 29.145 ;
        RECT 210.005 28.945 210.325 29.005 ;
        RECT 211.400 28.960 211.690 29.005 ;
        RECT 171.840 28.620 172.130 28.850 ;
        RECT 171.915 28.465 172.055 28.620 ;
        RECT 174.585 28.605 174.905 28.865 ;
        RECT 175.520 28.805 175.810 28.850 ;
        RECT 178.725 28.805 179.045 28.865 ;
        RECT 175.520 28.665 179.045 28.805 ;
        RECT 175.520 28.620 175.810 28.665 ;
        RECT 178.725 28.605 179.045 28.665 ;
        RECT 180.580 28.620 180.870 28.850 ;
        RECT 185.165 28.805 185.485 28.865 ;
        RECT 186.560 28.805 186.850 28.850 ;
        RECT 185.165 28.665 186.850 28.805 ;
        RECT 172.300 28.465 172.590 28.510 ;
        RECT 171.915 28.325 172.590 28.465 ;
        RECT 180.655 28.465 180.795 28.620 ;
        RECT 185.165 28.605 185.485 28.665 ;
        RECT 186.560 28.620 186.850 28.665 ;
        RECT 191.605 28.605 191.925 28.865 ;
        RECT 200.345 28.805 200.665 28.865 ;
        RECT 204.040 28.805 204.330 28.850 ;
        RECT 200.345 28.665 204.330 28.805 ;
        RECT 200.345 28.605 200.665 28.665 ;
        RECT 204.040 28.620 204.330 28.665 ;
        RECT 183.800 28.465 184.090 28.510 ;
        RECT 180.655 28.325 184.090 28.465 ;
        RECT 172.300 28.280 172.590 28.325 ;
        RECT 183.800 28.280 184.090 28.325 ;
        RECT 199.540 28.465 199.830 28.510 ;
        RECT 202.660 28.465 202.950 28.510 ;
        RECT 204.550 28.465 204.840 28.510 ;
        RECT 199.540 28.325 204.840 28.465 ;
        RECT 199.540 28.280 199.830 28.325 ;
        RECT 202.660 28.280 202.950 28.325 ;
        RECT 204.550 28.280 204.840 28.325 ;
        RECT 164.005 27.925 164.325 28.185 ;
        RECT 188.400 28.125 188.690 28.170 ;
        RECT 189.305 28.125 189.625 28.185 ;
        RECT 188.400 27.985 189.625 28.125 ;
        RECT 188.400 27.940 188.690 27.985 ;
        RECT 189.305 27.925 189.625 27.985 ;
        RECT 162.095 27.305 311.135 27.785 ;
        RECT 170.905 27.105 171.225 27.165 ;
        RECT 171.380 27.105 171.670 27.150 ;
        RECT 170.905 26.965 171.670 27.105 ;
        RECT 170.905 26.905 171.225 26.965 ;
        RECT 171.380 26.920 171.670 26.965 ;
        RECT 174.585 27.105 174.905 27.165 ;
        RECT 175.520 27.105 175.810 27.150 ;
        RECT 174.585 26.965 175.810 27.105 ;
        RECT 174.585 26.905 174.905 26.965 ;
        RECT 175.520 26.920 175.810 26.965 ;
        RECT 189.765 27.105 190.085 27.165 ;
        RECT 192.540 27.105 192.830 27.150 ;
        RECT 189.765 26.965 192.830 27.105 ;
        RECT 189.765 26.905 190.085 26.965 ;
        RECT 192.540 26.920 192.830 26.965 ;
        RECT 198.505 26.905 198.825 27.165 ;
        RECT 208.640 27.105 208.930 27.150 ;
        RECT 212.305 27.105 212.625 27.165 ;
        RECT 208.640 26.965 212.625 27.105 ;
        RECT 208.640 26.920 208.930 26.965 ;
        RECT 212.305 26.905 212.625 26.965 ;
        RECT 186.545 26.765 186.865 26.825 ;
        RECT 198.595 26.765 198.735 26.905 ;
        RECT 186.545 26.625 198.735 26.765 ;
        RECT 186.545 26.565 186.865 26.625 ;
        RECT 174.600 26.425 174.890 26.470 ;
        RECT 175.505 26.425 175.825 26.485 ;
        RECT 174.600 26.285 175.825 26.425 ;
        RECT 174.600 26.240 174.890 26.285 ;
        RECT 175.505 26.225 175.825 26.285 ;
        RECT 176.885 26.425 177.205 26.485 ;
        RECT 178.280 26.425 178.570 26.470 ;
        RECT 176.885 26.285 178.570 26.425 ;
        RECT 176.885 26.225 177.205 26.285 ;
        RECT 178.280 26.240 178.570 26.285 ;
        RECT 189.305 26.225 189.625 26.485 ;
        RECT 205.880 26.425 206.170 26.470 ;
        RECT 206.785 26.425 207.105 26.485 ;
        RECT 205.880 26.285 207.105 26.425 ;
        RECT 205.880 26.240 206.170 26.285 ;
        RECT 206.785 26.225 207.105 26.285 ;
        RECT 199.885 25.885 200.205 26.145 ;
        RECT 162.095 24.585 311.135 25.065 ;
        RECT 162.095 21.865 311.135 22.345 ;
        RECT 162.095 19.145 311.135 19.625 ;
        RECT 135.120 14.050 138.400 18.845 ;
        RECT 146.290 14.050 155.900 18.845 ;
        RECT 162.095 16.425 311.135 16.905 ;
        RECT 135.120 4.900 155.900 14.050 ;
        RECT 162.095 13.705 311.135 14.185 ;
        RECT 4.100 4.100 155.900 4.900 ;
      LAYER met2 ;
        RECT 45.340 224.760 45.740 225.560 ;
        RECT 64.710 225.410 217.040 225.710 ;
        RECT 64.710 225.310 65.510 225.410 ;
        RECT 59.190 224.760 59.990 225.160 ;
        RECT 67.470 224.810 207.380 225.110 ;
        RECT 67.470 224.710 68.270 224.810 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.210 197.720 224.510 ;
        RECT 70.230 224.110 71.030 224.210 ;
        RECT 72.990 223.610 188.060 223.910 ;
        RECT 72.990 223.510 73.790 223.610 ;
        RECT 75.700 223.010 178.400 223.310 ;
        RECT 75.700 222.910 76.500 223.010 ;
        RECT 78.545 222.410 168.740 222.710 ;
        RECT 78.545 222.310 79.345 222.410 ;
        RECT 83.980 221.810 164.500 222.110 ;
        RECT 83.980 221.710 84.780 221.810 ;
        RECT 86.740 221.210 163.500 221.510 ;
        RECT 164.100 221.310 164.500 221.810 ;
        RECT 86.740 221.110 87.540 221.210 ;
        RECT 92.260 220.610 162.500 220.910 ;
        RECT 163.100 220.710 163.500 221.210 ;
        RECT 92.260 220.510 93.060 220.610 ;
        RECT 162.100 220.110 162.500 220.610 ;
        RECT 6.200 211.890 7.800 215.090 ;
        RECT 9.570 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 9.495 208.765 51.905 210.765 ;
        RECT 9.495 205.765 45.165 207.765 ;
        RECT 51.315 207.460 51.905 208.765 ;
        RECT 9.495 202.765 48.270 204.765 ;
        RECT 9.495 198.745 48.270 200.745 ;
        RECT 9.495 195.745 45.165 197.745 ;
        RECT 9.495 192.745 46.670 194.745 ;
        RECT 9.495 187.420 15.245 188.980 ;
        RECT 16.515 188.295 45.165 190.295 ;
        RECT 52.860 188.465 54.245 190.570 ;
        RECT 16.515 184.775 56.920 186.775 ;
        RECT 6.200 180.050 7.800 183.250 ;
        RECT 9.495 182.570 15.245 184.130 ;
        RECT 16.515 181.255 46.670 183.255 ;
        RECT 5.910 176.050 7.510 179.250 ;
        RECT 57.020 178.865 57.820 178.990 ;
        RECT 9.500 177.365 58.420 178.865 ;
        RECT 53.870 176.720 54.670 176.890 ;
        RECT 9.500 175.220 54.670 176.720 ;
        RECT 9.500 172.820 54.670 174.320 ;
        RECT 53.870 172.640 54.670 172.820 ;
        RECT 52.220 171.920 53.020 172.040 ;
        RECT 9.500 170.420 53.020 171.920 ;
        RECT 63.470 170.855 65.220 217.105 ;
        RECT 66.220 170.855 67.970 217.105 ;
        RECT 68.970 170.855 70.720 217.105 ;
        RECT 71.720 170.855 73.470 217.105 ;
        RECT 74.470 170.855 76.220 217.105 ;
        RECT 77.220 170.855 78.970 217.105 ;
        RECT 79.970 170.115 81.970 217.845 ;
        RECT 106.340 217.515 107.940 219.915 ;
        RECT 109.240 219.705 111.675 220.105 ;
        RECT 113.270 219.705 115.705 220.105 ;
        RECT 117.300 219.705 119.735 220.105 ;
        RECT 121.330 219.705 123.765 220.105 ;
        RECT 125.360 219.705 127.795 220.105 ;
        RECT 129.390 219.705 131.825 220.105 ;
        RECT 133.420 219.705 135.855 220.105 ;
        RECT 137.450 219.705 139.885 220.105 ;
        RECT 141.480 219.705 143.915 220.105 ;
        RECT 145.510 219.705 147.945 220.105 ;
        RECT 149.540 219.705 151.975 220.105 ;
        RECT 109.240 217.705 109.640 219.705 ;
        RECT 110.530 217.705 110.930 219.305 ;
        RECT 111.820 217.295 112.220 219.305 ;
        RECT 113.270 217.705 113.670 219.705 ;
        RECT 114.560 217.705 114.960 219.305 ;
        RECT 115.850 217.295 116.250 219.305 ;
        RECT 117.300 217.705 117.700 219.705 ;
        RECT 118.590 217.705 118.990 219.305 ;
        RECT 119.880 217.295 120.280 219.305 ;
        RECT 121.330 217.705 121.730 219.705 ;
        RECT 122.620 217.705 123.020 219.305 ;
        RECT 123.910 217.295 124.310 219.305 ;
        RECT 125.360 217.705 125.760 219.705 ;
        RECT 126.650 217.705 127.050 219.305 ;
        RECT 127.940 217.295 128.340 219.305 ;
        RECT 129.390 217.705 129.790 219.705 ;
        RECT 130.680 217.705 131.080 219.305 ;
        RECT 131.970 217.295 132.370 219.305 ;
        RECT 133.420 217.705 133.820 219.705 ;
        RECT 134.710 217.705 135.110 219.305 ;
        RECT 136.000 217.295 136.400 219.305 ;
        RECT 137.450 217.705 137.850 219.705 ;
        RECT 138.740 217.705 139.140 219.305 ;
        RECT 140.030 217.295 140.430 219.305 ;
        RECT 141.480 217.705 141.880 219.705 ;
        RECT 142.770 217.705 143.170 219.305 ;
        RECT 144.060 217.295 144.460 219.305 ;
        RECT 145.510 217.705 145.910 219.705 ;
        RECT 146.800 217.705 147.200 219.305 ;
        RECT 148.090 217.295 148.490 219.305 ;
        RECT 149.540 217.705 149.940 219.705 ;
        RECT 150.830 217.705 151.230 219.305 ;
        RECT 152.120 217.295 152.520 219.305 ;
        RECT 82.970 170.855 84.720 217.105 ;
        RECT 85.720 170.855 87.470 217.105 ;
        RECT 88.470 170.855 90.220 217.105 ;
        RECT 91.220 170.855 92.970 217.105 ;
        RECT 93.970 170.855 95.720 217.105 ;
        RECT 96.720 170.855 98.470 217.105 ;
        RECT 109.785 216.895 112.220 217.295 ;
        RECT 113.815 216.895 116.250 217.295 ;
        RECT 117.845 216.895 120.280 217.295 ;
        RECT 121.875 216.895 124.310 217.295 ;
        RECT 125.905 216.895 128.340 217.295 ;
        RECT 129.935 216.895 132.370 217.295 ;
        RECT 133.965 216.895 136.400 217.295 ;
        RECT 137.995 216.895 140.430 217.295 ;
        RECT 142.025 216.895 144.460 217.295 ;
        RECT 146.055 216.895 148.490 217.295 ;
        RECT 150.085 216.895 152.520 217.295 ;
        RECT 106.415 210.540 108.015 213.740 ;
        RECT 110.530 209.640 110.930 211.240 ;
        RECT 114.560 209.640 114.960 211.240 ;
        RECT 118.590 209.640 118.990 211.240 ;
        RECT 122.620 209.640 123.020 211.240 ;
        RECT 126.650 209.640 127.050 211.240 ;
        RECT 130.680 209.640 131.080 211.240 ;
        RECT 134.710 209.640 135.110 211.240 ;
        RECT 138.740 209.640 139.140 211.240 ;
        RECT 142.770 209.640 143.170 211.240 ;
        RECT 146.800 209.640 147.200 211.240 ;
        RECT 150.830 209.640 151.230 211.240 ;
        RECT 111.820 205.955 112.220 206.755 ;
        RECT 115.850 205.955 116.250 206.755 ;
        RECT 119.880 205.955 120.280 206.755 ;
        RECT 123.910 205.955 124.310 206.755 ;
        RECT 127.940 205.955 128.340 206.755 ;
        RECT 131.970 205.955 132.370 206.755 ;
        RECT 136.000 205.955 136.400 206.755 ;
        RECT 140.030 205.955 140.430 206.755 ;
        RECT 144.060 205.955 144.460 206.755 ;
        RECT 148.090 205.955 148.490 206.755 ;
        RECT 152.120 205.955 152.520 206.755 ;
        RECT 109.240 204.745 111.675 205.545 ;
        RECT 113.270 204.745 115.705 205.545 ;
        RECT 117.300 204.745 119.735 205.545 ;
        RECT 121.330 204.745 123.765 205.545 ;
        RECT 125.360 204.745 127.795 205.545 ;
        RECT 129.390 204.745 131.825 205.545 ;
        RECT 133.420 204.745 135.855 205.545 ;
        RECT 137.450 204.745 139.885 205.545 ;
        RECT 141.480 204.745 143.915 205.545 ;
        RECT 145.510 204.745 147.945 205.545 ;
        RECT 149.540 204.745 151.975 205.545 ;
        RECT 108.540 202.425 108.940 202.625 ;
        RECT 109.785 202.425 110.385 204.345 ;
        RECT 108.540 202.025 110.385 202.425 ;
        RECT 108.540 201.825 108.940 202.025 ;
        RECT 109.785 199.970 110.385 202.025 ;
        RECT 111.075 199.970 111.675 204.745 ;
        RECT 112.570 202.425 112.970 202.625 ;
        RECT 113.815 202.425 114.415 204.345 ;
        RECT 112.570 202.025 114.415 202.425 ;
        RECT 112.570 201.825 112.970 202.025 ;
        RECT 113.815 199.970 114.415 202.025 ;
        RECT 115.105 199.970 115.705 204.745 ;
        RECT 116.600 202.425 117.000 202.625 ;
        RECT 117.845 202.425 118.445 204.345 ;
        RECT 116.600 202.025 118.445 202.425 ;
        RECT 116.600 201.825 117.000 202.025 ;
        RECT 117.845 199.970 118.445 202.025 ;
        RECT 119.135 199.970 119.735 204.745 ;
        RECT 120.630 202.425 121.030 202.625 ;
        RECT 121.875 202.425 122.475 204.345 ;
        RECT 120.630 202.025 122.475 202.425 ;
        RECT 120.630 201.825 121.030 202.025 ;
        RECT 121.875 199.970 122.475 202.025 ;
        RECT 123.165 199.970 123.765 204.745 ;
        RECT 124.660 202.425 125.060 202.625 ;
        RECT 125.905 202.425 126.505 204.345 ;
        RECT 124.660 202.025 126.505 202.425 ;
        RECT 124.660 201.825 125.060 202.025 ;
        RECT 125.905 199.970 126.505 202.025 ;
        RECT 127.195 199.970 127.795 204.745 ;
        RECT 128.690 202.425 129.090 202.625 ;
        RECT 129.935 202.425 130.535 204.345 ;
        RECT 128.690 202.025 130.535 202.425 ;
        RECT 128.690 201.825 129.090 202.025 ;
        RECT 129.935 199.970 130.535 202.025 ;
        RECT 131.225 199.970 131.825 204.745 ;
        RECT 132.720 202.425 133.120 202.625 ;
        RECT 133.965 202.425 134.565 204.345 ;
        RECT 132.720 202.025 134.565 202.425 ;
        RECT 132.720 201.825 133.120 202.025 ;
        RECT 133.965 199.970 134.565 202.025 ;
        RECT 135.255 199.970 135.855 204.745 ;
        RECT 136.750 202.425 137.150 202.625 ;
        RECT 137.995 202.425 138.595 204.345 ;
        RECT 136.750 202.025 138.595 202.425 ;
        RECT 136.750 201.825 137.150 202.025 ;
        RECT 137.995 199.970 138.595 202.025 ;
        RECT 139.285 199.970 139.885 204.745 ;
        RECT 140.780 202.425 141.180 202.625 ;
        RECT 142.025 202.425 142.625 204.345 ;
        RECT 140.780 202.025 142.625 202.425 ;
        RECT 140.780 201.825 141.180 202.025 ;
        RECT 142.025 199.970 142.625 202.025 ;
        RECT 143.315 199.970 143.915 204.745 ;
        RECT 144.810 202.425 145.210 202.625 ;
        RECT 146.055 202.425 146.655 204.345 ;
        RECT 144.810 202.025 146.655 202.425 ;
        RECT 144.810 201.825 145.210 202.025 ;
        RECT 146.055 199.970 146.655 202.025 ;
        RECT 147.345 199.970 147.945 204.745 ;
        RECT 148.840 202.425 149.240 202.625 ;
        RECT 150.085 202.425 150.685 204.345 ;
        RECT 148.840 202.025 150.685 202.425 ;
        RECT 148.840 201.825 149.240 202.025 ;
        RECT 150.085 199.970 150.685 202.025 ;
        RECT 151.375 199.970 151.975 204.745 ;
        RECT 168.460 202.290 168.740 222.410 ;
        RECT 178.120 202.290 178.400 223.010 ;
        RECT 187.780 202.290 188.060 223.610 ;
        RECT 197.440 202.290 197.720 224.210 ;
        RECT 207.100 202.290 207.380 224.810 ;
        RECT 216.760 202.290 217.040 225.410 ;
        RECT 246.615 225.060 247.015 225.660 ;
        RECT 226.420 224.460 226.700 224.510 ;
        RECT 236.020 224.460 236.420 225.060 ;
        RECT 226.360 223.860 226.760 224.460 ;
        RECT 226.420 202.290 226.700 223.860 ;
        RECT 236.080 202.290 236.360 224.460 ;
        RECT 246.665 218.450 246.965 225.060 ;
        RECT 246.615 217.650 247.015 218.450 ;
        RECT 168.530 201.140 168.670 202.290 ;
        RECT 178.190 201.140 178.330 202.290 ;
        RECT 180.700 201.305 182.240 201.675 ;
        RECT 187.850 201.140 187.990 202.290 ;
        RECT 197.510 201.140 197.650 202.290 ;
        RECT 207.170 201.140 207.310 202.290 ;
        RECT 216.830 201.140 216.970 202.290 ;
        RECT 226.490 201.140 226.630 202.290 ;
        RECT 236.150 201.140 236.290 202.290 ;
        RECT 168.470 200.820 168.730 201.140 ;
        RECT 178.130 200.820 178.390 201.140 ;
        RECT 187.790 200.820 188.050 201.140 ;
        RECT 197.450 200.820 197.710 201.140 ;
        RECT 207.110 200.820 207.370 201.140 ;
        RECT 216.770 200.820 217.030 201.140 ;
        RECT 226.430 200.820 226.690 201.140 ;
        RECT 236.090 200.820 236.350 201.140 ;
        RECT 166.630 199.800 166.890 200.120 ;
        RECT 170.310 199.800 170.570 200.120 ;
        RECT 178.590 199.800 178.850 200.120 ;
        RECT 191.470 199.800 191.730 200.120 ;
        RECT 197.910 199.800 198.170 200.120 ;
        RECT 208.950 199.800 209.210 200.120 ;
        RECT 217.230 199.800 217.490 200.120 ;
        RECT 226.890 199.800 227.150 200.120 ;
        RECT 236.090 199.800 236.350 200.120 ;
        RECT 109.240 194.440 109.640 199.685 ;
        RECT 109.240 194.040 110.255 194.440 ;
        RECT 109.240 191.285 109.640 192.885 ;
        RECT 110.530 187.540 110.930 198.905 ;
        RECT 111.820 194.440 112.220 199.685 ;
        RECT 111.205 194.040 112.220 194.440 ;
        RECT 113.270 194.440 113.670 199.685 ;
        RECT 113.270 194.040 114.285 194.440 ;
        RECT 111.820 191.285 112.220 192.885 ;
        RECT 113.270 191.285 113.670 192.885 ;
        RECT 114.560 187.540 114.960 198.905 ;
        RECT 115.850 194.440 116.250 199.685 ;
        RECT 115.235 194.040 116.250 194.440 ;
        RECT 117.300 194.440 117.700 199.685 ;
        RECT 117.300 194.040 118.315 194.440 ;
        RECT 115.850 191.285 116.250 192.885 ;
        RECT 117.300 191.285 117.700 192.885 ;
        RECT 118.590 187.540 118.990 198.905 ;
        RECT 119.880 194.440 120.280 199.685 ;
        RECT 119.265 194.040 120.280 194.440 ;
        RECT 121.330 194.440 121.730 199.685 ;
        RECT 121.330 194.040 122.345 194.440 ;
        RECT 119.880 191.285 120.280 192.885 ;
        RECT 121.330 191.285 121.730 192.885 ;
        RECT 122.620 187.540 123.020 198.905 ;
        RECT 123.910 194.440 124.310 199.685 ;
        RECT 123.295 194.040 124.310 194.440 ;
        RECT 125.360 194.440 125.760 199.685 ;
        RECT 125.360 194.040 126.375 194.440 ;
        RECT 123.910 191.285 124.310 192.885 ;
        RECT 125.360 191.285 125.760 192.885 ;
        RECT 126.650 187.540 127.050 198.905 ;
        RECT 127.940 194.440 128.340 199.685 ;
        RECT 127.325 194.040 128.340 194.440 ;
        RECT 129.390 194.440 129.790 199.685 ;
        RECT 129.390 194.040 130.405 194.440 ;
        RECT 127.940 191.285 128.340 192.885 ;
        RECT 129.390 191.285 129.790 192.885 ;
        RECT 130.680 187.540 131.080 198.905 ;
        RECT 131.970 194.440 132.370 199.685 ;
        RECT 131.355 194.040 132.370 194.440 ;
        RECT 133.420 194.440 133.820 199.685 ;
        RECT 133.420 194.040 134.435 194.440 ;
        RECT 131.970 191.285 132.370 192.885 ;
        RECT 133.420 191.285 133.820 192.885 ;
        RECT 134.710 187.540 135.110 198.905 ;
        RECT 136.000 194.440 136.400 199.685 ;
        RECT 135.385 194.040 136.400 194.440 ;
        RECT 137.450 194.440 137.850 199.685 ;
        RECT 137.450 194.040 138.465 194.440 ;
        RECT 136.000 191.285 136.400 192.885 ;
        RECT 137.450 191.285 137.850 192.885 ;
        RECT 138.740 187.540 139.140 198.905 ;
        RECT 140.030 194.440 140.430 199.685 ;
        RECT 139.415 194.040 140.430 194.440 ;
        RECT 141.480 194.440 141.880 199.685 ;
        RECT 141.480 194.040 142.495 194.440 ;
        RECT 140.030 191.285 140.430 192.885 ;
        RECT 141.480 191.285 141.880 192.885 ;
        RECT 142.770 187.540 143.170 198.905 ;
        RECT 144.060 194.440 144.460 199.685 ;
        RECT 143.445 194.040 144.460 194.440 ;
        RECT 145.510 194.440 145.910 199.685 ;
        RECT 145.510 194.040 146.525 194.440 ;
        RECT 144.060 191.285 144.460 192.885 ;
        RECT 145.510 191.285 145.910 192.885 ;
        RECT 146.800 187.540 147.200 198.905 ;
        RECT 148.090 194.440 148.490 199.685 ;
        RECT 147.475 194.040 148.490 194.440 ;
        RECT 149.540 194.440 149.940 199.685 ;
        RECT 149.540 194.040 150.555 194.440 ;
        RECT 148.090 191.285 148.490 192.885 ;
        RECT 149.540 191.285 149.940 192.885 ;
        RECT 150.830 187.540 151.230 198.905 ;
        RECT 152.120 194.440 152.520 199.685 ;
        RECT 166.690 197.935 166.830 199.800 ;
        RECT 166.620 197.565 166.900 197.935 ;
        RECT 151.505 194.040 152.520 194.440 ;
        RECT 152.120 191.285 152.520 192.885 ;
        RECT 167.540 192.805 167.820 193.175 ;
        RECT 167.610 190.260 167.750 192.805 ;
        RECT 170.370 190.260 170.510 199.800 ;
        RECT 174.450 199.120 174.710 199.440 ;
        RECT 174.510 192.495 174.650 199.120 ;
        RECT 178.650 192.980 178.790 199.800 ;
        RECT 184.000 198.585 185.540 198.955 ;
        RECT 180.700 195.865 182.240 196.235 ;
        RECT 181.350 193.680 181.610 194.000 ;
        RECT 178.590 192.660 178.850 192.980 ;
        RECT 173.530 191.980 173.790 192.300 ;
        RECT 174.440 192.125 174.720 192.495 ;
        RECT 173.070 190.960 173.330 191.280 ;
        RECT 167.550 189.940 167.810 190.260 ;
        RECT 170.310 189.940 170.570 190.260 ;
        RECT 171.690 189.260 171.950 189.580 ;
        RECT 166.630 188.920 166.890 189.240 ;
        RECT 161.590 188.380 162.390 188.430 ;
        RECT 166.690 188.415 166.830 188.920 ;
        RECT 158.335 188.080 162.390 188.380 ;
        RECT 109.240 184.370 109.640 184.770 ;
        RECT 153.565 184.765 155.165 187.965 ;
        RECT 158.335 187.580 158.735 188.080 ;
        RECT 161.590 188.030 162.390 188.080 ;
        RECT 166.620 188.045 166.900 188.415 ;
        RECT 168.000 187.365 168.280 187.735 ;
        RECT 168.010 187.220 168.270 187.365 ;
        RECT 168.470 187.220 168.730 187.540 ;
        RECT 167.550 186.200 167.810 186.520 ;
        RECT 167.610 184.820 167.750 186.200 ;
        RECT 167.550 184.500 167.810 184.820 ;
        RECT 109.240 183.970 154.345 184.370 ;
        RECT 153.945 183.570 154.345 183.970 ;
        RECT 168.530 183.800 168.670 187.220 ;
        RECT 168.930 186.540 169.190 186.860 ;
        RECT 170.310 186.540 170.570 186.860 ;
        RECT 168.990 184.820 169.130 186.540 ;
        RECT 169.850 185.750 170.110 185.840 ;
        RECT 169.450 185.610 170.110 185.750 ;
        RECT 168.930 184.500 169.190 184.820 ;
        RECT 166.630 183.480 166.890 183.800 ;
        RECT 168.470 183.480 168.730 183.800 ;
        RECT 166.690 179.040 166.830 183.480 ;
        RECT 167.090 181.100 167.350 181.420 ;
        RECT 161.590 178.860 162.390 178.910 ;
        RECT 157.560 178.560 162.390 178.860 ;
        RECT 166.630 178.720 166.890 179.040 ;
        RECT 167.150 178.895 167.290 181.100 ;
        RECT 168.990 180.255 169.130 184.500 ;
        RECT 169.450 181.615 169.590 185.610 ;
        RECT 169.850 185.520 170.110 185.610 ;
        RECT 169.850 183.480 170.110 183.800 ;
        RECT 169.910 182.100 170.050 183.480 ;
        RECT 169.850 181.780 170.110 182.100 ;
        RECT 169.380 181.245 169.660 181.615 ;
        RECT 169.390 180.650 169.650 180.740 ;
        RECT 170.370 180.650 170.510 186.540 ;
        RECT 170.770 185.520 171.030 185.840 ;
        RECT 170.830 181.420 170.970 185.520 ;
        RECT 171.750 184.220 171.890 189.260 ;
        RECT 172.150 188.920 172.410 189.240 ;
        RECT 172.210 184.820 172.350 188.920 ;
        RECT 172.610 188.240 172.870 188.560 ;
        RECT 172.150 184.500 172.410 184.820 ;
        RECT 171.750 184.080 172.350 184.220 ;
        RECT 171.230 183.140 171.490 183.460 ;
        RECT 171.690 183.140 171.950 183.460 ;
        RECT 170.770 181.100 171.030 181.420 ;
        RECT 169.390 180.510 170.510 180.650 ;
        RECT 169.390 180.420 169.650 180.510 ;
        RECT 168.920 179.885 169.200 180.255 ;
        RECT 169.450 178.895 169.590 180.420 ;
        RECT 115.265 175.815 117.965 176.215 ;
        RECT 119.885 175.815 122.585 176.215 ;
        RECT 124.505 175.815 127.205 176.215 ;
        RECT 129.125 175.815 131.825 176.215 ;
        RECT 133.745 175.815 136.445 176.215 ;
        RECT 138.365 175.815 141.065 176.215 ;
        RECT 142.985 175.815 145.685 176.215 ;
        RECT 147.605 175.815 150.305 176.215 ;
        RECT 151.155 175.010 152.755 178.210 ;
        RECT 157.560 178.060 157.960 178.560 ;
        RECT 161.590 178.510 162.390 178.560 ;
        RECT 167.080 178.525 167.360 178.895 ;
        RECT 169.380 178.525 169.660 178.895 ;
        RECT 170.830 178.360 170.970 181.100 ;
        RECT 171.290 179.380 171.430 183.140 ;
        RECT 171.750 182.100 171.890 183.140 ;
        RECT 171.690 181.780 171.950 182.100 ;
        RECT 172.210 180.935 172.350 184.080 ;
        RECT 172.140 180.565 172.420 180.935 ;
        RECT 171.230 179.060 171.490 179.380 ;
        RECT 172.670 178.360 172.810 188.240 ;
        RECT 173.130 182.100 173.270 190.960 ;
        RECT 173.070 181.780 173.330 182.100 ;
        RECT 173.590 181.500 173.730 191.980 ;
        RECT 173.990 189.600 174.250 189.920 ;
        RECT 173.130 181.360 173.730 181.500 ;
        RECT 168.470 178.040 168.730 178.360 ;
        RECT 170.770 178.040 171.030 178.360 ;
        RECT 172.150 178.040 172.410 178.360 ;
        RECT 172.610 178.040 172.870 178.360 ;
        RECT 168.530 176.855 168.670 178.040 ;
        RECT 172.210 177.680 172.350 178.040 ;
        RECT 172.150 177.360 172.410 177.680 ;
        RECT 168.460 176.485 168.740 176.855 ;
        RECT 173.130 176.290 173.270 181.360 ;
        RECT 174.050 176.290 174.190 189.600 ;
        RECT 174.510 183.800 174.650 192.125 ;
        RECT 175.370 191.980 175.630 192.300 ;
        RECT 177.670 191.980 177.930 192.300 ;
        RECT 178.590 191.980 178.850 192.300 ;
        RECT 179.050 191.980 179.310 192.300 ;
        RECT 180.890 192.210 181.150 192.300 ;
        RECT 179.570 192.070 181.150 192.210 ;
        RECT 174.910 190.960 175.170 191.280 ;
        RECT 174.970 189.240 175.110 190.960 ;
        RECT 174.910 188.920 175.170 189.240 ;
        RECT 175.430 188.160 175.570 191.980 ;
        RECT 175.830 191.300 176.090 191.620 ;
        RECT 174.970 188.020 175.570 188.160 ;
        RECT 174.450 183.480 174.710 183.800 ;
        RECT 174.450 180.080 174.710 180.400 ;
        RECT 174.510 178.360 174.650 180.080 ;
        RECT 174.450 178.040 174.710 178.360 ;
        RECT 174.970 176.290 175.110 188.020 ;
        RECT 175.890 186.860 176.030 191.300 ;
        RECT 177.730 191.280 177.870 191.980 ;
        RECT 178.130 191.300 178.390 191.620 ;
        RECT 177.670 190.960 177.930 191.280 ;
        RECT 176.290 188.920 176.550 189.240 ;
        RECT 176.350 187.540 176.490 188.920 ;
        RECT 177.670 188.580 177.930 188.900 ;
        RECT 176.290 187.220 176.550 187.540 ;
        RECT 175.830 186.540 176.090 186.860 ;
        RECT 175.370 183.480 175.630 183.800 ;
        RECT 175.890 183.655 176.030 186.540 ;
        RECT 176.350 184.480 176.490 187.220 ;
        RECT 177.730 186.860 177.870 188.580 ;
        RECT 178.190 188.560 178.330 191.300 ;
        RECT 178.130 188.240 178.390 188.560 ;
        RECT 177.670 186.540 177.930 186.860 ;
        RECT 176.750 185.520 177.010 185.840 ;
        RECT 176.290 184.160 176.550 184.480 ;
        RECT 175.430 180.400 175.570 183.480 ;
        RECT 175.820 183.285 176.100 183.655 ;
        RECT 176.290 183.480 176.550 183.800 ;
        RECT 175.820 182.605 176.100 182.975 ;
        RECT 175.890 182.100 176.030 182.605 ;
        RECT 175.830 181.780 176.090 182.100 ;
        RECT 175.820 181.245 176.100 181.615 ;
        RECT 175.370 180.080 175.630 180.400 ;
        RECT 175.360 179.205 175.640 179.575 ;
        RECT 175.370 179.060 175.630 179.205 ;
        RECT 175.890 176.290 176.030 181.245 ;
        RECT 176.350 179.380 176.490 183.480 ;
        RECT 176.810 182.975 176.950 185.520 ;
        RECT 177.200 183.965 177.480 184.335 ;
        RECT 177.270 183.800 177.410 183.965 ;
        RECT 177.730 183.800 177.870 186.540 ;
        RECT 178.130 185.860 178.390 186.180 ;
        RECT 178.190 184.140 178.330 185.860 ;
        RECT 178.650 184.820 178.790 191.980 ;
        RECT 179.110 191.815 179.250 191.980 ;
        RECT 179.040 191.445 179.320 191.815 ;
        RECT 179.110 189.580 179.250 191.445 ;
        RECT 179.050 189.260 179.310 189.580 ;
        RECT 179.040 188.725 179.320 189.095 ;
        RECT 178.590 184.500 178.850 184.820 ;
        RECT 178.130 183.820 178.390 184.140 ;
        RECT 177.210 183.480 177.470 183.800 ;
        RECT 177.670 183.480 177.930 183.800 ;
        RECT 176.740 182.605 177.020 182.975 ;
        RECT 176.750 181.780 177.010 182.100 ;
        RECT 176.290 179.060 176.550 179.380 ;
        RECT 176.810 176.290 176.950 181.780 ;
        RECT 177.210 181.100 177.470 181.420 ;
        RECT 177.270 176.320 177.410 181.100 ;
        RECT 177.730 181.080 177.870 183.480 ;
        RECT 178.130 183.140 178.390 183.460 ;
        RECT 177.670 180.760 177.930 181.080 ;
        RECT 177.670 180.080 177.930 180.400 ;
        RECT 177.730 179.575 177.870 180.080 ;
        RECT 177.660 179.205 177.940 179.575 ;
        RECT 177.670 178.720 177.930 179.040 ;
        RECT 114.835 172.120 118.395 174.820 ;
        RECT 119.155 172.120 123.015 174.820 ;
        RECT 123.775 172.120 127.635 174.820 ;
        RECT 128.395 172.120 132.255 174.820 ;
        RECT 133.015 172.120 136.875 174.820 ;
        RECT 137.635 172.120 141.495 174.820 ;
        RECT 142.255 172.120 146.115 174.820 ;
        RECT 146.875 172.120 150.735 174.820 ;
        RECT 57.020 169.775 57.820 169.890 ;
        RECT 9.500 168.275 58.420 169.775 ;
        RECT 9.500 165.715 56.920 166.715 ;
        RECT 103.350 164.990 103.750 170.890 ;
        RECT 105.930 168.490 106.330 170.890 ;
        RECT 9.500 163.915 55.070 164.915 ;
        RECT 102.625 164.590 103.750 164.990 ;
        RECT 104.640 164.790 105.040 167.190 ;
        RECT 107.380 164.990 107.780 170.890 ;
        RECT 109.960 168.490 110.360 170.890 ;
        RECT 115.625 169.795 117.605 170.845 ;
        RECT 119.155 169.795 119.755 172.120 ;
        RECT 115.625 169.195 119.755 169.795 ;
        RECT 120.245 169.795 122.225 170.845 ;
        RECT 123.775 169.795 124.375 172.120 ;
        RECT 120.245 169.195 124.375 169.795 ;
        RECT 124.865 169.795 126.845 170.845 ;
        RECT 128.395 169.795 128.995 172.120 ;
        RECT 124.865 169.195 128.995 169.795 ;
        RECT 129.485 169.795 131.465 170.845 ;
        RECT 133.015 169.795 133.615 172.120 ;
        RECT 129.485 169.195 133.615 169.795 ;
        RECT 134.105 169.795 136.085 170.845 ;
        RECT 137.635 169.795 138.235 172.120 ;
        RECT 134.105 169.195 138.235 169.795 ;
        RECT 138.725 169.795 140.705 170.845 ;
        RECT 142.255 169.795 142.855 172.120 ;
        RECT 138.725 169.195 142.855 169.795 ;
        RECT 143.345 169.795 145.325 170.845 ;
        RECT 146.875 169.795 147.475 172.120 ;
        RECT 143.345 169.195 147.475 169.795 ;
        RECT 115.625 168.145 117.605 169.195 ;
        RECT 120.245 168.145 122.225 169.195 ;
        RECT 124.865 168.145 126.845 169.195 ;
        RECT 129.485 168.145 131.465 169.195 ;
        RECT 134.105 168.145 136.085 169.195 ;
        RECT 138.725 168.145 140.705 169.195 ;
        RECT 143.345 168.145 145.325 169.195 ;
        RECT 147.965 168.145 150.345 170.845 ;
        RECT 106.655 164.590 107.780 164.990 ;
        RECT 108.670 164.790 109.070 167.190 ;
        RECT 9.500 162.115 51.610 163.115 ;
        RECT 9.500 159.815 53.170 161.315 ;
        RECT 2.705 157.015 51.610 159.015 ;
        RECT 2.705 1.285 3.505 157.015 ;
        RECT 9.500 154.715 53.170 156.215 ;
        RECT 9.500 152.915 51.610 153.915 ;
        RECT 9.500 151.115 55.070 152.115 ;
        RECT 74.940 151.875 86.100 155.595 ;
        RECT 9.500 149.315 56.520 150.315 ;
        RECT 51.580 145.090 53.180 148.290 ;
        RECT 71.585 145.090 73.185 148.290 ;
        RECT 74.940 148.155 78.660 151.875 ;
        RECT 80.100 149.595 80.930 150.425 ;
        RECT 82.380 148.155 86.100 151.875 ;
        RECT 102.625 149.850 103.025 164.590 ;
        RECT 103.350 162.940 104.365 163.340 ;
        RECT 105.315 162.940 106.330 163.340 ;
        RECT 103.350 159.695 103.750 162.940 ;
        RECT 105.930 160.395 106.330 162.940 ;
        RECT 104.190 159.795 106.330 160.395 ;
        RECT 104.190 159.410 104.495 159.795 ;
        RECT 105.930 159.695 106.330 159.795 ;
        RECT 103.895 154.535 104.495 159.410 ;
        RECT 105.185 155.035 105.785 159.410 ;
        RECT 103.895 153.935 106.330 154.535 ;
        RECT 103.350 150.640 103.750 153.565 ;
        RECT 105.930 152.190 106.330 153.935 ;
        RECT 103.895 151.790 106.330 152.190 ;
        RECT 103.895 151.015 104.495 151.790 ;
        RECT 105.185 150.640 105.785 151.415 ;
        RECT 103.350 150.240 105.785 150.640 ;
        RECT 106.655 149.850 107.055 164.590 ;
        RECT 107.380 162.940 108.395 163.340 ;
        RECT 109.345 162.940 110.360 163.340 ;
        RECT 107.380 159.695 107.780 162.940 ;
        RECT 109.960 160.395 110.360 162.940 ;
        RECT 108.220 159.795 110.360 160.395 ;
        RECT 108.220 159.410 108.525 159.795 ;
        RECT 109.960 159.695 110.360 159.795 ;
        RECT 107.925 154.535 108.525 159.410 ;
        RECT 109.215 155.035 109.815 159.410 ;
        RECT 107.925 153.935 110.360 154.535 ;
        RECT 107.380 150.640 107.780 153.565 ;
        RECT 109.960 152.190 110.360 153.935 ;
        RECT 107.925 151.790 110.360 152.190 ;
        RECT 107.925 151.015 108.525 151.790 ;
        RECT 109.215 150.640 109.815 151.415 ;
        RECT 107.380 150.240 109.815 150.640 ;
        RECT 102.625 149.450 103.750 149.850 ;
        RECT 74.940 144.435 86.100 148.155 ;
        RECT 20.350 141.375 20.750 142.975 ;
        RECT 11.195 139.800 23.015 140.200 ;
        RECT 11.195 137.185 11.795 139.800 ;
        RECT 14.860 138.370 21.050 138.770 ;
        RECT 14.860 137.585 15.260 138.370 ;
        RECT 20.650 137.970 21.050 138.370 ;
        RECT 14.130 137.185 16.020 137.585 ;
        RECT 16.805 137.185 18.955 137.585 ;
        RECT 16.805 136.875 17.205 137.185 ;
        RECT 11.940 136.275 15.275 136.875 ;
        RECT 16.165 136.275 17.205 136.875 ;
        RECT 5.910 132.225 7.510 135.425 ;
        RECT 13.485 133.130 14.085 135.875 ;
        RECT 13.385 132.330 14.185 133.130 ;
        RECT 16.805 129.110 17.205 136.275 ;
        RECT 19.100 136.125 20.750 136.725 ;
        RECT 16.805 128.710 17.605 129.110 ;
        RECT 19.100 128.925 19.500 136.125 ;
        RECT 22.615 134.120 23.015 139.800 ;
        RECT 24.255 135.155 25.755 143.745 ;
        RECT 27.765 135.155 29.265 143.745 ;
        RECT 36.055 135.155 37.555 143.745 ;
        RECT 44.345 135.155 45.845 143.745 ;
        RECT 52.635 135.155 54.135 143.745 ;
        RECT 56.145 135.155 57.645 143.745 ;
        RECT 103.350 143.435 103.750 149.450 ;
        RECT 104.640 147.135 105.040 149.535 ;
        RECT 106.655 149.450 107.780 149.850 ;
        RECT 105.930 143.435 106.330 145.835 ;
        RECT 107.380 143.435 107.780 149.450 ;
        RECT 108.670 147.135 109.070 149.535 ;
        RECT 109.960 143.435 110.360 145.835 ;
        RECT 116.310 143.410 116.910 168.145 ;
        RECT 120.930 147.550 121.530 168.145 ;
        RECT 125.550 159.440 126.150 168.145 ;
        RECT 125.550 158.840 128.940 159.440 ;
        RECT 120.930 146.950 126.935 147.550 ;
        RECT 122.645 144.030 124.245 144.830 ;
        RECT 128.340 144.540 128.940 158.840 ;
        RECT 130.170 148.610 130.770 168.145 ;
        RECT 134.795 164.330 135.395 168.145 ;
        RECT 133.685 163.140 134.485 163.740 ;
        RECT 133.785 155.610 134.385 163.140 ;
        RECT 136.775 161.650 137.575 162.450 ;
        RECT 134.695 159.460 135.495 160.260 ;
        RECT 139.410 157.075 140.010 168.145 ;
        RECT 144.035 163.040 144.635 168.145 ;
        RECT 146.855 164.430 147.655 165.030 ;
        RECT 143.935 161.650 144.735 162.450 ;
        RECT 145.525 159.460 146.325 160.260 ;
        RECT 141.615 158.550 142.415 159.150 ;
        RECT 138.070 156.475 140.010 157.075 ;
        RECT 133.285 155.010 134.885 155.610 ;
        RECT 133.275 151.400 134.875 152.200 ;
        RECT 133.275 150.230 134.875 151.030 ;
        RECT 138.070 149.760 138.670 156.475 ;
        RECT 141.715 152.110 142.315 158.550 ;
        RECT 141.215 151.905 142.815 152.110 ;
        RECT 140.950 151.505 143.050 151.905 ;
        RECT 133.285 149.160 138.670 149.760 ;
        RECT 130.170 148.010 134.430 148.610 ;
        RECT 130.615 146.830 132.215 147.630 ;
        RECT 133.285 147.410 134.885 148.010 ;
        RECT 138.525 147.310 140.125 148.110 ;
        RECT 128.340 143.940 134.885 144.540 ;
        RECT 138.525 143.820 140.125 144.620 ;
        RECT 116.310 142.810 132.215 143.410 ;
        RECT 141.215 143.240 142.815 144.040 ;
        RECT 141.215 141.990 142.815 142.790 ;
        RECT 146.955 142.730 147.555 164.430 ;
        RECT 148.655 158.450 149.255 168.145 ;
        RECT 146.455 142.640 148.055 142.730 ;
        RECT 146.195 142.240 148.295 142.640 ;
        RECT 146.455 142.130 148.055 142.240 ;
        RECT 104.640 139.365 152.360 140.165 ;
        RECT 97.200 137.420 147.750 138.220 ;
        RECT 107.380 135.525 132.465 136.325 ;
        RECT 22.615 133.320 23.415 134.120 ;
        RECT 56.145 133.555 77.110 135.155 ;
        RECT 80.120 133.320 137.265 134.120 ;
        RECT 137.945 133.410 144.375 133.810 ;
        RECT 21.615 131.745 135.665 132.545 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 142.980 131.990 143.630 132.590 ;
        RECT 27.065 129.995 134.065 130.795 ;
        RECT 19.100 128.125 101.315 128.925 ;
        RECT 6.200 124.285 7.800 127.485 ;
        RECT 65.865 124.285 67.465 127.485 ;
        RECT 121.565 124.285 123.165 127.485 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 141.700 125.690 142.100 127.290 ;
        RECT 142.980 126.815 143.230 131.990 ;
        RECT 144.025 131.050 144.375 133.410 ;
        RECT 143.725 129.545 144.425 131.050 ;
        RECT 153.945 129.545 154.345 129.945 ;
        RECT 143.725 129.145 154.345 129.545 ;
        RECT 143.725 127.640 144.425 129.145 ;
        RECT 142.980 126.215 143.630 126.815 ;
        RECT 10.025 122.800 70.175 123.810 ;
        RECT 71.775 122.750 114.165 123.850 ;
        RECT 10.025 120.300 70.175 122.300 ;
        RECT 71.775 121.250 114.165 122.350 ;
        RECT 115.905 121.575 128.935 123.145 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 10.025 117.800 70.175 119.800 ;
        RECT 71.775 119.750 114.165 120.850 ;
        RECT 71.775 118.250 114.165 119.350 ;
        RECT 10.025 115.300 70.175 117.300 ;
        RECT 71.775 116.750 114.165 117.850 ;
        RECT 115.905 117.075 128.935 118.645 ;
        RECT 141.900 116.370 150.745 117.170 ;
        RECT 71.775 115.250 114.165 116.350 ;
        RECT 10.025 112.780 70.175 114.800 ;
        RECT 71.775 112.730 114.165 114.850 ;
        RECT 136.465 114.770 144.870 115.570 ;
        RECT 173.060 115.285 173.340 176.290 ;
        RECT 115.905 112.615 128.935 114.185 ;
        RECT 10.025 110.280 70.175 112.280 ;
        RECT 71.775 111.230 114.165 112.330 ;
        RECT 133.265 111.795 141.675 112.595 ;
        RECT 10.025 107.780 70.175 109.780 ;
        RECT 71.775 109.730 114.165 110.830 ;
        RECT 140.875 110.315 141.675 111.795 ;
        RECT 144.070 110.315 144.870 114.770 ;
        RECT 164.025 115.005 173.340 115.285 ;
        RECT 71.775 108.230 114.165 109.330 ;
        RECT 115.905 108.115 128.935 109.685 ;
        RECT 139.560 109.515 142.995 110.315 ;
        RECT 136.295 108.925 138.400 109.515 ;
        RECT 10.025 105.280 70.175 107.280 ;
        RECT 71.775 106.730 114.165 107.830 ;
        RECT 71.775 105.230 114.165 106.330 ;
        RECT 10.025 103.770 70.175 104.780 ;
        RECT 71.775 103.730 114.165 104.830 ;
        RECT 115.905 103.655 128.935 105.225 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 10.025 91.525 128.935 92.775 ;
        RECT 10.025 89.640 128.935 91.140 ;
        RECT 10.025 85.640 128.935 88.640 ;
        RECT 136.295 86.115 138.400 90.215 ;
        RECT 10.025 83.140 128.935 84.640 ;
        RECT 10.025 81.505 128.935 82.755 ;
        RECT 10.025 79.620 128.935 81.120 ;
        RECT 136.295 80.265 138.400 85.535 ;
        RECT 139.560 82.025 140.860 109.515 ;
        RECT 141.695 91.385 142.995 109.515 ;
        RECT 141.290 90.795 143.395 91.385 ;
        RECT 139.155 81.435 141.260 82.025 ;
        RECT 10.025 75.620 128.935 78.620 ;
        RECT 136.295 75.585 138.400 79.685 ;
        RECT 10.025 73.120 128.935 74.620 ;
        RECT 10.025 71.485 128.935 72.735 ;
        RECT 10.025 69.600 128.935 71.100 ;
        RECT 136.295 70.905 138.400 75.005 ;
        RECT 10.025 65.600 128.935 68.600 ;
        RECT 136.295 66.225 138.400 70.325 ;
        RECT 10.025 63.100 128.935 64.600 ;
        RECT 10.025 61.465 128.935 62.715 ;
        RECT 10.025 59.580 128.935 61.080 ;
        RECT 136.295 60.375 138.400 65.645 ;
        RECT 10.025 55.580 128.935 58.580 ;
        RECT 136.295 55.695 138.400 59.795 ;
        RECT 10.025 53.080 128.935 54.580 ;
        RECT 10.025 51.445 128.935 52.695 ;
        RECT 136.295 51.015 138.400 55.115 ;
        RECT 12.915 45.565 14.515 47.165 ;
        RECT 90.715 45.565 92.315 47.165 ;
        RECT 136.295 46.335 138.400 50.435 ;
        RECT 6.200 41.635 7.800 44.835 ;
        RECT 136.295 40.485 138.400 45.755 ;
        RECT 143.835 42.245 145.135 110.315 ;
        RECT 164.025 109.225 164.305 115.005 ;
        RECT 173.980 114.705 174.260 176.290 ;
        RECT 166.325 114.425 174.260 114.705 ;
        RECT 166.325 109.225 166.605 114.425 ;
        RECT 174.900 114.125 175.180 176.290 ;
        RECT 168.625 113.845 175.180 114.125 ;
        RECT 168.625 109.225 168.905 113.845 ;
        RECT 175.820 113.545 176.100 176.290 ;
        RECT 170.925 113.265 176.100 113.545 ;
        RECT 170.925 109.225 171.205 113.265 ;
        RECT 176.740 112.965 177.020 176.290 ;
        RECT 177.210 176.000 177.470 176.320 ;
        RECT 177.730 176.290 177.870 178.720 ;
        RECT 173.225 112.685 177.020 112.965 ;
        RECT 173.225 109.225 173.505 112.685 ;
        RECT 177.660 112.385 177.940 176.290 ;
        RECT 178.190 175.980 178.330 183.140 ;
        RECT 178.590 181.440 178.850 181.760 ;
        RECT 178.650 179.380 178.790 181.440 ;
        RECT 179.110 181.420 179.250 188.725 ;
        RECT 179.050 181.100 179.310 181.420 ;
        RECT 179.050 180.420 179.310 180.740 ;
        RECT 179.110 180.255 179.250 180.420 ;
        RECT 179.040 179.885 179.320 180.255 ;
        RECT 178.590 179.060 178.850 179.380 ;
        RECT 178.580 178.525 178.860 178.895 ;
        RECT 178.650 176.290 178.790 178.525 ;
        RECT 179.570 176.290 179.710 192.070 ;
        RECT 180.890 191.980 181.150 192.070 ;
        RECT 181.410 191.280 181.550 193.680 ;
        RECT 181.800 192.805 182.080 193.175 ;
        RECT 184.000 193.145 185.540 193.515 ;
        RECT 191.530 192.980 191.670 199.800 ;
        RECT 197.970 192.980 198.110 199.800 ;
        RECT 207.570 193.680 207.830 194.000 ;
        RECT 181.870 192.640 182.010 192.805 ;
        RECT 182.270 192.660 182.530 192.980 ;
        RECT 191.470 192.660 191.730 192.980 ;
        RECT 197.910 192.660 198.170 192.980 ;
        RECT 181.810 192.320 182.070 192.640 ;
        RECT 181.810 191.870 182.070 191.960 ;
        RECT 182.330 191.870 182.470 192.660 ;
        RECT 184.100 192.210 184.380 192.495 ;
        RECT 188.250 192.320 188.510 192.640 ;
        RECT 184.100 192.125 185.230 192.210 ;
        RECT 184.110 192.070 185.230 192.125 ;
        RECT 184.110 191.980 184.370 192.070 ;
        RECT 181.810 191.730 182.470 191.870 ;
        RECT 181.810 191.640 182.070 191.730 ;
        RECT 182.730 191.640 182.990 191.960 ;
        RECT 181.350 190.960 181.610 191.280 ;
        RECT 180.700 190.425 182.240 190.795 ;
        RECT 179.970 188.920 180.230 189.240 ;
        RECT 180.890 188.920 181.150 189.240 ;
        RECT 182.270 189.150 182.530 189.240 ;
        RECT 182.790 189.150 182.930 191.640 ;
        RECT 183.190 190.960 183.450 191.280 ;
        RECT 183.250 190.340 183.390 190.960 ;
        RECT 183.250 190.200 184.310 190.340 ;
        RECT 182.270 189.010 182.930 189.150 ;
        RECT 182.270 188.920 182.530 189.010 ;
        RECT 180.030 187.735 180.170 188.920 ;
        RECT 179.960 187.365 180.240 187.735 ;
        RECT 180.950 187.540 181.090 188.920 ;
        RECT 182.270 188.240 182.530 188.560 ;
        RECT 184.170 188.470 184.310 190.200 ;
        RECT 185.090 189.580 185.230 192.070 ;
        RECT 185.950 191.980 186.210 192.300 ;
        RECT 186.010 189.920 186.150 191.980 ;
        RECT 185.950 189.600 186.210 189.920 ;
        RECT 185.030 189.490 185.290 189.580 ;
        RECT 185.030 189.350 185.690 189.490 ;
        RECT 185.030 189.260 185.290 189.350 ;
        RECT 185.020 188.725 185.300 189.095 ;
        RECT 185.090 188.560 185.230 188.725 ;
        RECT 183.250 188.330 184.310 188.470 ;
        RECT 182.330 187.540 182.470 188.240 ;
        RECT 180.890 187.220 181.150 187.540 ;
        RECT 182.270 187.220 182.530 187.540 ;
        RECT 179.970 186.880 180.230 187.200 ;
        RECT 180.430 187.055 180.690 187.200 ;
        RECT 180.030 182.100 180.170 186.880 ;
        RECT 180.420 186.685 180.700 187.055 ;
        RECT 180.950 186.860 181.090 187.220 ;
        RECT 180.890 186.540 181.150 186.860 ;
        RECT 182.270 186.540 182.530 186.860 ;
        RECT 182.330 185.750 182.470 186.540 ;
        RECT 182.330 185.610 182.930 185.750 ;
        RECT 180.700 184.985 182.240 185.355 ;
        RECT 180.890 183.480 181.150 183.800 ;
        RECT 180.430 182.800 180.690 183.120 ;
        RECT 179.970 181.780 180.230 182.100 ;
        RECT 180.490 180.740 180.630 182.800 ;
        RECT 180.950 181.420 181.090 183.480 ;
        RECT 181.340 183.285 181.620 183.655 ;
        RECT 182.270 183.480 182.530 183.800 ;
        RECT 181.410 181.760 181.550 183.285 ;
        RECT 181.810 183.140 182.070 183.460 ;
        RECT 181.350 181.440 181.610 181.760 ;
        RECT 181.870 181.420 182.010 183.140 ;
        RECT 182.330 181.615 182.470 183.480 ;
        RECT 180.890 181.100 181.150 181.420 ;
        RECT 181.810 181.100 182.070 181.420 ;
        RECT 182.260 181.245 182.540 181.615 ;
        RECT 180.430 180.420 180.690 180.740 ;
        RECT 180.700 179.545 182.240 179.915 ;
        RECT 180.430 178.380 180.690 178.700 ;
        RECT 181.340 178.525 181.620 178.895 ;
        RECT 182.790 178.780 182.930 185.610 ;
        RECT 183.250 181.420 183.390 188.330 ;
        RECT 185.030 188.240 185.290 188.560 ;
        RECT 185.550 188.470 185.690 189.350 ;
        RECT 186.410 188.920 186.670 189.240 ;
        RECT 186.870 188.920 187.130 189.240 ;
        RECT 185.550 188.330 186.150 188.470 ;
        RECT 184.000 187.705 185.540 188.075 ;
        RECT 186.010 187.450 186.150 188.330 ;
        RECT 186.470 187.540 186.610 188.920 ;
        RECT 185.550 187.310 186.150 187.450 ;
        RECT 184.570 186.880 184.830 187.200 ;
        RECT 183.650 186.540 183.910 186.860 ;
        RECT 183.190 181.100 183.450 181.420 ;
        RECT 183.710 180.820 183.850 186.540 ;
        RECT 184.110 185.520 184.370 185.840 ;
        RECT 184.170 183.800 184.310 185.520 ;
        RECT 184.630 183.800 184.770 186.880 ;
        RECT 185.030 186.540 185.290 186.860 ;
        RECT 185.090 184.335 185.230 186.540 ;
        RECT 185.020 183.965 185.300 184.335 ;
        RECT 184.110 183.480 184.370 183.800 ;
        RECT 184.570 183.480 184.830 183.800 ;
        RECT 185.550 183.460 185.690 187.310 ;
        RECT 186.410 187.220 186.670 187.540 ;
        RECT 186.930 187.200 187.070 188.920 ;
        RECT 187.330 188.240 187.590 188.560 ;
        RECT 186.870 186.880 187.130 187.200 ;
        RECT 185.950 186.540 186.210 186.860 ;
        RECT 185.490 183.140 185.750 183.460 ;
        RECT 184.000 182.265 185.540 182.635 ;
        RECT 185.490 181.100 185.750 181.420 ;
        RECT 182.330 178.640 182.930 178.780 ;
        RECT 183.250 180.680 183.850 180.820 ;
        RECT 179.970 178.040 180.230 178.360 ;
        RECT 178.130 175.660 178.390 175.980 ;
        RECT 175.525 112.105 177.940 112.385 ;
        RECT 175.525 109.225 175.805 112.105 ;
        RECT 178.580 111.805 178.860 176.290 ;
        RECT 177.825 111.525 178.860 111.805 ;
        RECT 179.500 111.805 179.780 176.290 ;
        RECT 180.030 175.640 180.170 178.040 ;
        RECT 180.490 176.290 180.630 178.380 ;
        RECT 181.410 178.360 181.550 178.525 ;
        RECT 181.350 178.040 181.610 178.360 ;
        RECT 180.890 177.360 181.150 177.680 ;
        RECT 181.810 177.360 182.070 177.680 ;
        RECT 179.970 175.320 180.230 175.640 ;
        RECT 180.420 112.385 180.700 176.290 ;
        RECT 180.950 174.960 181.090 177.360 ;
        RECT 181.340 176.485 181.620 176.855 ;
        RECT 181.410 176.290 181.550 176.485 ;
        RECT 180.890 174.640 181.150 174.960 ;
        RECT 181.340 112.965 181.620 176.290 ;
        RECT 181.870 175.300 182.010 177.360 ;
        RECT 182.330 176.290 182.470 178.640 ;
        RECT 182.730 177.700 182.990 178.020 ;
        RECT 182.790 176.855 182.930 177.700 ;
        RECT 182.720 176.485 183.000 176.855 ;
        RECT 183.250 176.290 183.390 180.680 ;
        RECT 184.570 180.255 184.830 180.400 ;
        RECT 183.640 179.885 183.920 180.255 ;
        RECT 184.560 179.885 184.840 180.255 ;
        RECT 183.710 176.570 183.850 179.885 ;
        RECT 185.550 179.575 185.690 181.100 ;
        RECT 185.480 179.205 185.760 179.575 ;
        RECT 184.000 176.825 185.540 177.195 ;
        RECT 185.490 176.570 185.750 176.660 ;
        RECT 183.710 176.430 184.310 176.570 ;
        RECT 184.170 176.290 184.310 176.430 ;
        RECT 185.090 176.430 185.750 176.570 ;
        RECT 185.090 176.290 185.230 176.430 ;
        RECT 185.490 176.340 185.750 176.430 ;
        RECT 186.010 176.290 186.150 186.540 ;
        RECT 187.390 186.375 187.530 188.240 ;
        RECT 187.790 186.540 188.050 186.860 ;
        RECT 187.320 186.005 187.600 186.375 ;
        RECT 186.410 185.520 186.670 185.840 ;
        RECT 187.330 185.520 187.590 185.840 ;
        RECT 186.470 183.800 186.610 185.520 ;
        RECT 186.870 184.500 187.130 184.820 ;
        RECT 186.930 184.335 187.070 184.500 ;
        RECT 186.860 183.965 187.140 184.335 ;
        RECT 186.410 183.480 186.670 183.800 ;
        RECT 186.875 183.480 187.135 183.800 ;
        RECT 186.930 182.975 187.070 183.480 ;
        RECT 186.860 182.605 187.140 182.975 ;
        RECT 186.400 181.925 186.680 182.295 ;
        RECT 186.410 181.780 186.670 181.925 ;
        RECT 186.860 181.245 187.140 181.615 ;
        RECT 186.410 178.040 186.670 178.360 ;
        RECT 181.810 174.980 182.070 175.300 ;
        RECT 182.260 113.545 182.540 176.290 ;
        RECT 183.180 114.125 183.460 176.290 ;
        RECT 184.100 114.705 184.380 176.290 ;
        RECT 185.020 115.285 185.300 176.290 ;
        RECT 185.940 115.865 186.220 176.290 ;
        RECT 186.470 175.980 186.610 178.040 ;
        RECT 186.930 176.290 187.070 181.245 ;
        RECT 187.390 178.360 187.530 185.520 ;
        RECT 187.330 178.040 187.590 178.360 ;
        RECT 187.330 177.360 187.590 177.680 ;
        RECT 187.390 176.320 187.530 177.360 ;
        RECT 186.410 175.660 186.670 175.980 ;
        RECT 186.860 116.445 187.140 176.290 ;
        RECT 187.330 176.000 187.590 176.320 ;
        RECT 187.850 176.290 187.990 186.540 ;
        RECT 188.310 182.100 188.450 192.320 ;
        RECT 194.230 191.980 194.490 192.300 ;
        RECT 198.830 191.980 199.090 192.300 ;
        RECT 193.770 191.815 194.030 191.960 ;
        RECT 193.760 191.445 194.040 191.815 ;
        RECT 194.290 191.190 194.430 191.980 ;
        RECT 193.830 191.050 194.430 191.190 ;
        RECT 189.170 188.920 189.430 189.240 ;
        RECT 190.090 189.150 190.350 189.240 ;
        RECT 189.690 189.010 190.350 189.150 ;
        RECT 189.230 187.540 189.370 188.920 ;
        RECT 189.170 187.220 189.430 187.540 ;
        RECT 189.690 187.200 189.830 189.010 ;
        RECT 190.090 188.920 190.350 189.010 ;
        RECT 191.010 189.150 191.270 189.240 ;
        RECT 191.010 189.010 193.510 189.150 ;
        RECT 191.010 188.920 191.270 189.010 ;
        RECT 189.630 186.880 189.890 187.200 ;
        RECT 189.170 186.540 189.430 186.860 ;
        RECT 188.710 185.520 188.970 185.840 ;
        RECT 188.770 182.100 188.910 185.520 ;
        RECT 188.250 181.780 188.510 182.100 ;
        RECT 188.710 181.780 188.970 182.100 ;
        RECT 188.250 181.100 188.510 181.420 ;
        RECT 188.310 178.700 188.450 181.100 ;
        RECT 189.230 180.820 189.370 186.540 ;
        RECT 189.690 183.800 189.830 186.880 ;
        RECT 190.090 186.540 190.350 186.860 ;
        RECT 191.470 186.540 191.730 186.860 ;
        RECT 190.150 185.695 190.290 186.540 ;
        RECT 190.080 185.325 190.360 185.695 ;
        RECT 191.000 183.965 191.280 184.335 ;
        RECT 189.630 183.655 189.890 183.800 ;
        RECT 189.620 183.285 189.900 183.655 ;
        RECT 190.090 183.140 190.350 183.460 ;
        RECT 188.770 180.680 189.370 180.820 ;
        RECT 188.250 178.380 188.510 178.700 ;
        RECT 188.770 176.290 188.910 180.680 ;
        RECT 190.150 179.380 190.290 183.140 ;
        RECT 191.070 183.120 191.210 183.965 ;
        RECT 191.010 182.800 191.270 183.120 ;
        RECT 190.540 181.245 190.820 181.615 ;
        RECT 190.550 181.100 190.810 181.245 ;
        RECT 191.010 181.100 191.270 181.420 ;
        RECT 191.070 180.740 191.210 181.100 ;
        RECT 191.010 180.420 191.270 180.740 ;
        RECT 190.090 179.060 190.350 179.380 ;
        RECT 191.010 178.040 191.270 178.360 ;
        RECT 190.090 177.700 190.350 178.020 ;
        RECT 189.620 177.165 189.900 177.535 ;
        RECT 189.690 176.290 189.830 177.165 ;
        RECT 187.780 117.025 188.060 176.290 ;
        RECT 188.700 117.605 188.980 176.290 ;
        RECT 189.620 118.185 189.900 176.290 ;
        RECT 190.150 174.620 190.290 177.700 ;
        RECT 191.070 177.535 191.210 178.040 ;
        RECT 191.000 177.165 191.280 177.535 ;
        RECT 190.610 176.430 191.210 176.570 ;
        RECT 190.610 176.290 190.750 176.430 ;
        RECT 190.090 174.300 190.350 174.620 ;
        RECT 190.540 118.765 190.820 176.290 ;
        RECT 191.070 176.175 191.210 176.430 ;
        RECT 191.530 176.290 191.670 186.540 ;
        RECT 192.390 186.200 192.650 186.520 ;
        RECT 191.930 184.160 192.190 184.480 ;
        RECT 191.990 180.400 192.130 184.160 ;
        RECT 192.450 184.140 192.590 186.200 ;
        RECT 192.850 185.520 193.110 185.840 ;
        RECT 192.390 183.820 192.650 184.140 ;
        RECT 192.380 182.605 192.660 182.975 ;
        RECT 192.450 182.100 192.590 182.605 ;
        RECT 192.390 181.780 192.650 182.100 ;
        RECT 191.930 180.080 192.190 180.400 ;
        RECT 192.380 178.525 192.660 178.895 ;
        RECT 191.930 178.040 192.190 178.360 ;
        RECT 191.990 176.660 192.130 178.040 ;
        RECT 192.450 177.420 192.590 178.525 ;
        RECT 192.910 178.360 193.050 185.520 ;
        RECT 193.370 184.820 193.510 189.010 ;
        RECT 193.830 187.540 193.970 191.050 ;
        RECT 198.890 190.260 199.030 191.980 ;
        RECT 200.210 191.640 200.470 191.960 ;
        RECT 198.830 189.940 199.090 190.260 ;
        RECT 196.520 189.405 196.800 189.775 ;
        RECT 200.270 189.580 200.410 191.640 ;
        RECT 206.650 191.300 206.910 191.620 ;
        RECT 202.970 190.960 203.230 191.280 ;
        RECT 196.590 189.240 196.730 189.405 ;
        RECT 200.210 189.260 200.470 189.580 ;
        RECT 196.530 188.920 196.790 189.240 ;
        RECT 194.230 188.580 194.490 188.900 ;
        RECT 193.770 187.220 194.030 187.540 ;
        RECT 193.830 186.860 193.970 187.220 ;
        RECT 193.770 186.540 194.030 186.860 ;
        RECT 193.830 186.180 193.970 186.540 ;
        RECT 193.770 185.860 194.030 186.180 ;
        RECT 193.310 184.500 193.570 184.820 ;
        RECT 193.830 183.800 193.970 185.860 ;
        RECT 194.290 184.140 194.430 188.580 ;
        RECT 199.750 188.240 200.010 188.560 ;
        RECT 199.810 187.200 199.950 188.240 ;
        RECT 199.750 186.880 200.010 187.200 ;
        RECT 195.150 186.540 195.410 186.860 ;
        RECT 196.070 186.540 196.330 186.860 ;
        RECT 198.370 186.770 198.630 186.860 ;
        RECT 197.970 186.630 198.630 186.770 ;
        RECT 194.230 183.820 194.490 184.140 ;
        RECT 193.770 183.480 194.030 183.800 ;
        RECT 193.770 183.030 194.030 183.120 ;
        RECT 193.370 182.890 194.030 183.030 ;
        RECT 192.850 178.040 193.110 178.360 ;
        RECT 193.370 178.270 193.510 182.890 ;
        RECT 193.770 182.800 194.030 182.890 ;
        RECT 194.290 181.080 194.430 183.820 ;
        RECT 194.690 182.800 194.950 183.120 ;
        RECT 194.230 180.760 194.490 181.080 ;
        RECT 193.760 179.205 194.040 179.575 ;
        RECT 194.290 179.380 194.430 180.760 ;
        RECT 193.830 178.610 193.970 179.205 ;
        RECT 194.230 179.060 194.490 179.380 ;
        RECT 194.750 179.040 194.890 182.800 ;
        RECT 195.210 182.100 195.350 186.540 ;
        RECT 195.610 182.800 195.870 183.120 ;
        RECT 195.150 181.780 195.410 182.100 ;
        RECT 195.670 180.400 195.810 182.800 ;
        RECT 195.610 180.080 195.870 180.400 ;
        RECT 196.130 180.255 196.270 186.540 ;
        RECT 196.990 186.200 197.250 186.520 ;
        RECT 197.050 183.540 197.190 186.200 ;
        RECT 197.450 184.500 197.710 184.820 ;
        RECT 196.590 183.460 197.190 183.540 ;
        RECT 196.530 183.400 197.190 183.460 ;
        RECT 196.530 183.140 196.790 183.400 ;
        RECT 196.530 181.100 196.790 181.420 ;
        RECT 196.060 179.885 196.340 180.255 ;
        RECT 194.690 178.720 194.950 179.040 ;
        RECT 193.830 178.470 194.430 178.610 ;
        RECT 193.370 178.130 193.970 178.270 ;
        RECT 192.450 177.280 193.510 177.420 ;
        RECT 191.930 176.340 192.190 176.660 ;
        RECT 192.450 176.600 193.050 176.740 ;
        RECT 192.450 176.290 192.590 176.600 ;
        RECT 191.000 175.805 191.280 176.175 ;
        RECT 191.460 119.345 191.740 176.290 ;
        RECT 192.380 119.925 192.660 176.290 ;
        RECT 192.910 175.640 193.050 176.600 ;
        RECT 193.370 176.290 193.510 177.280 ;
        RECT 192.850 175.320 193.110 175.640 ;
        RECT 193.300 120.505 193.580 176.290 ;
        RECT 193.830 174.960 193.970 178.130 ;
        RECT 194.290 176.290 194.430 178.470 ;
        RECT 194.750 176.430 195.350 176.570 ;
        RECT 193.770 174.640 194.030 174.960 ;
        RECT 194.220 121.085 194.500 176.290 ;
        RECT 194.750 174.620 194.890 176.430 ;
        RECT 195.210 176.290 195.350 176.430 ;
        RECT 195.670 176.430 196.270 176.570 ;
        RECT 194.690 174.300 194.950 174.620 ;
        RECT 195.140 121.665 195.420 176.290 ;
        RECT 195.670 175.980 195.810 176.430 ;
        RECT 196.130 176.290 196.270 176.430 ;
        RECT 195.610 175.660 195.870 175.980 ;
        RECT 196.060 122.245 196.340 176.290 ;
        RECT 196.590 175.300 196.730 181.100 ;
        RECT 197.510 180.820 197.650 184.500 ;
        RECT 197.970 183.800 198.110 186.630 ;
        RECT 198.370 186.540 198.630 186.630 ;
        RECT 199.290 186.540 199.550 186.860 ;
        RECT 200.200 186.685 200.480 187.055 ;
        RECT 201.120 186.685 201.400 187.055 ;
        RECT 200.210 186.540 200.470 186.685 ;
        RECT 198.830 185.860 199.090 186.180 ;
        RECT 197.910 183.480 198.170 183.800 ;
        RECT 198.370 183.140 198.630 183.460 ;
        RECT 198.430 182.100 198.570 183.140 ;
        RECT 198.370 181.780 198.630 182.100 ;
        RECT 198.890 181.615 199.030 185.860 ;
        RECT 198.820 181.245 199.100 181.615 ;
        RECT 197.050 180.680 197.650 180.820 ;
        RECT 197.910 180.760 198.170 181.080 ;
        RECT 197.050 176.290 197.190 180.680 ;
        RECT 197.970 179.380 198.110 180.760 ;
        RECT 199.350 179.380 199.490 186.540 ;
        RECT 201.190 184.480 201.330 186.685 ;
        RECT 202.510 186.540 202.770 186.860 ;
        RECT 202.570 184.820 202.710 186.540 ;
        RECT 202.510 184.500 202.770 184.820 ;
        RECT 201.130 184.160 201.390 184.480 ;
        RECT 200.670 183.480 200.930 183.800 ;
        RECT 199.750 182.800 200.010 183.120 ;
        RECT 197.910 179.060 198.170 179.380 ;
        RECT 199.290 179.060 199.550 179.380 ;
        RECT 197.900 177.165 198.180 177.535 ;
        RECT 197.970 176.290 198.110 177.165 ;
        RECT 198.370 176.570 198.630 176.660 ;
        RECT 198.370 176.430 199.030 176.570 ;
        RECT 198.370 176.340 198.630 176.430 ;
        RECT 198.890 176.290 199.030 176.430 ;
        RECT 199.810 176.290 199.950 182.800 ;
        RECT 200.200 181.925 200.480 182.295 ;
        RECT 200.210 181.780 200.470 181.925 ;
        RECT 200.730 176.290 200.870 183.480 ;
        RECT 201.130 182.800 201.390 183.120 ;
        RECT 201.590 182.800 201.850 183.120 ;
        RECT 201.190 181.760 201.330 182.800 ;
        RECT 201.130 181.440 201.390 181.760 ;
        RECT 201.130 178.380 201.390 178.700 ;
        RECT 201.190 178.215 201.330 178.380 ;
        RECT 201.650 178.360 201.790 182.800 ;
        RECT 202.510 181.100 202.770 181.420 ;
        RECT 202.050 180.760 202.310 181.080 ;
        RECT 202.110 178.700 202.250 180.760 ;
        RECT 202.050 178.380 202.310 178.700 ;
        RECT 201.120 177.845 201.400 178.215 ;
        RECT 201.590 178.040 201.850 178.360 ;
        RECT 201.590 177.360 201.850 177.680 ;
        RECT 201.650 176.290 201.790 177.360 ;
        RECT 196.530 174.980 196.790 175.300 ;
        RECT 196.980 122.825 197.260 176.290 ;
        RECT 197.900 123.405 198.180 176.290 ;
        RECT 198.820 123.985 199.100 176.290 ;
        RECT 199.740 124.565 200.020 176.290 ;
        RECT 200.660 125.145 200.940 176.290 ;
        RECT 201.580 125.725 201.860 176.290 ;
        RECT 202.110 175.980 202.250 178.380 ;
        RECT 202.570 176.290 202.710 181.100 ;
        RECT 203.030 178.895 203.170 190.960 ;
        RECT 203.430 182.800 203.690 183.120 ;
        RECT 203.490 179.380 203.630 182.800 ;
        RECT 206.190 181.440 206.450 181.760 ;
        RECT 205.270 181.100 205.530 181.420 ;
        RECT 203.430 179.060 203.690 179.380 ;
        RECT 202.960 178.525 203.240 178.895 ;
        RECT 203.430 178.040 203.690 178.360 ;
        RECT 204.350 178.040 204.610 178.360 ;
        RECT 203.490 176.290 203.630 178.040 ;
        RECT 204.410 176.290 204.550 178.040 ;
        RECT 205.330 176.290 205.470 181.100 ;
        RECT 206.250 176.290 206.390 181.440 ;
        RECT 206.710 179.380 206.850 191.300 ;
        RECT 207.110 185.860 207.370 186.180 ;
        RECT 207.170 181.080 207.310 185.860 ;
        RECT 207.110 180.760 207.370 181.080 ;
        RECT 206.650 179.060 206.910 179.380 ;
        RECT 207.630 178.700 207.770 193.680 ;
        RECT 209.010 187.540 209.150 199.800 ;
        RECT 216.770 192.320 217.030 192.640 ;
        RECT 210.330 189.260 210.590 189.580 ;
        RECT 208.950 187.220 209.210 187.540 ;
        RECT 209.410 187.220 209.670 187.540 ;
        RECT 209.470 185.840 209.610 187.220 ;
        RECT 210.390 186.860 210.530 189.260 ;
        RECT 210.790 188.920 211.050 189.240 ;
        RECT 210.850 187.200 210.990 188.920 ;
        RECT 210.790 186.880 211.050 187.200 ;
        RECT 211.250 186.880 211.510 187.200 ;
        RECT 210.330 186.540 210.590 186.860 ;
        RECT 209.870 186.375 210.130 186.520 ;
        RECT 209.860 186.005 210.140 186.375 ;
        RECT 211.310 186.090 211.450 186.880 ;
        RECT 213.090 186.540 213.350 186.860 ;
        RECT 215.390 186.540 215.650 186.860 ;
        RECT 212.170 186.200 212.430 186.520 ;
        RECT 212.630 186.200 212.890 186.520 ;
        RECT 210.850 185.950 211.450 186.090 ;
        RECT 209.410 185.520 209.670 185.840 ;
        RECT 209.870 185.520 210.130 185.840 ;
        RECT 209.410 183.820 209.670 184.140 ;
        RECT 208.490 183.710 208.750 183.800 ;
        RECT 208.490 183.570 209.150 183.710 ;
        RECT 208.490 183.480 208.750 183.570 ;
        RECT 207.570 178.380 207.830 178.700 ;
        RECT 207.170 176.660 207.770 176.740 ;
        RECT 207.170 176.600 207.830 176.660 ;
        RECT 207.170 176.290 207.310 176.600 ;
        RECT 207.570 176.340 207.830 176.600 ;
        RECT 208.090 176.600 208.690 176.740 ;
        RECT 208.090 176.290 208.230 176.600 ;
        RECT 208.550 176.320 208.690 176.600 ;
        RECT 202.050 175.660 202.310 175.980 ;
        RECT 202.500 126.305 202.780 176.290 ;
        RECT 203.420 126.885 203.700 176.290 ;
        RECT 204.340 127.465 204.620 176.290 ;
        RECT 205.260 128.045 205.540 176.290 ;
        RECT 206.180 128.625 206.460 176.290 ;
        RECT 207.100 129.205 207.380 176.290 ;
        RECT 208.020 129.785 208.300 176.290 ;
        RECT 208.490 176.000 208.750 176.320 ;
        RECT 209.010 176.290 209.150 183.570 ;
        RECT 209.470 180.740 209.610 183.820 ;
        RECT 209.410 180.420 209.670 180.740 ;
        RECT 209.470 179.380 209.610 180.420 ;
        RECT 209.410 179.060 209.670 179.380 ;
        RECT 209.930 176.290 210.070 185.520 ;
        RECT 210.850 182.860 210.990 185.950 ;
        RECT 211.710 185.520 211.970 185.840 ;
        RECT 211.250 184.730 211.510 184.820 ;
        RECT 211.770 184.730 211.910 185.520 ;
        RECT 211.250 184.590 211.910 184.730 ;
        RECT 211.250 184.500 211.510 184.590 ;
        RECT 211.710 183.820 211.970 184.140 ;
        RECT 211.770 182.975 211.910 183.820 ;
        RECT 210.850 182.720 211.450 182.860 ;
        RECT 210.330 181.780 210.590 182.100 ;
        RECT 210.780 181.925 211.060 182.295 ;
        RECT 210.390 181.615 210.530 181.780 ;
        RECT 210.320 181.245 210.600 181.615 ;
        RECT 210.330 178.380 210.590 178.700 ;
        RECT 210.390 178.215 210.530 178.380 ;
        RECT 210.320 177.845 210.600 178.215 ;
        RECT 210.850 176.290 210.990 181.925 ;
        RECT 211.310 177.590 211.450 182.720 ;
        RECT 211.700 182.605 211.980 182.975 ;
        RECT 211.700 181.925 211.980 182.295 ;
        RECT 211.770 181.080 211.910 181.925 ;
        RECT 212.230 181.080 212.370 186.200 ;
        RECT 211.710 180.760 211.970 181.080 ;
        RECT 212.170 180.760 212.430 181.080 ;
        RECT 212.160 179.205 212.440 179.575 ;
        RECT 211.710 178.270 211.970 178.360 ;
        RECT 212.230 178.270 212.370 179.205 ;
        RECT 211.710 178.130 212.370 178.270 ;
        RECT 211.710 178.040 211.970 178.130 ;
        RECT 211.310 177.450 211.910 177.590 ;
        RECT 211.770 176.290 211.910 177.450 ;
        RECT 212.690 176.290 212.830 186.200 ;
        RECT 213.150 185.695 213.290 186.540 ;
        RECT 213.080 185.325 213.360 185.695 ;
        RECT 214.930 185.520 215.190 185.840 ;
        RECT 213.090 184.500 213.350 184.820 ;
        RECT 213.150 184.140 213.290 184.500 ;
        RECT 214.990 184.140 215.130 185.520 ;
        RECT 213.090 183.820 213.350 184.140 ;
        RECT 214.010 184.050 214.270 184.140 ;
        RECT 214.010 183.910 214.670 184.050 ;
        RECT 214.010 183.820 214.270 183.910 ;
        RECT 213.090 180.990 213.350 181.080 ;
        RECT 214.530 180.990 214.670 183.910 ;
        RECT 214.930 183.820 215.190 184.140 ;
        RECT 213.090 180.850 214.670 180.990 ;
        RECT 213.090 180.760 213.350 180.850 ;
        RECT 213.150 178.215 213.290 180.760 ;
        RECT 214.000 179.885 214.280 180.255 ;
        RECT 213.550 179.290 213.810 179.380 ;
        RECT 214.070 179.290 214.210 179.885 ;
        RECT 213.550 179.150 214.210 179.290 ;
        RECT 214.460 179.205 214.740 179.575 ;
        RECT 213.550 179.060 213.810 179.150 ;
        RECT 214.530 178.610 214.670 179.205 ;
        RECT 214.930 179.060 215.190 179.380 ;
        RECT 214.990 178.700 215.130 179.060 ;
        RECT 214.070 178.470 214.670 178.610 ;
        RECT 214.070 178.270 214.210 178.470 ;
        RECT 214.930 178.380 215.190 178.700 ;
        RECT 213.080 177.845 213.360 178.215 ;
        RECT 213.610 178.130 214.210 178.270 ;
        RECT 213.610 176.290 213.750 178.130 ;
        RECT 215.450 178.100 215.590 186.540 ;
        RECT 216.830 184.820 216.970 192.320 ;
        RECT 217.290 190.260 217.430 199.800 ;
        RECT 225.970 190.960 226.230 191.280 ;
        RECT 226.030 190.260 226.170 190.960 ;
        RECT 226.950 190.260 227.090 199.800 ;
        RECT 232.410 190.960 232.670 191.280 ;
        RECT 217.230 189.940 217.490 190.260 ;
        RECT 225.970 189.940 226.230 190.260 ;
        RECT 226.890 189.940 227.150 190.260 ;
        RECT 225.050 189.660 225.310 189.920 ;
        RECT 224.650 189.600 225.310 189.660 ;
        RECT 231.490 189.600 231.750 189.920 ;
        RECT 224.650 189.520 225.250 189.600 ;
        RECT 218.150 186.880 218.410 187.200 ;
        RECT 219.990 186.880 220.250 187.200 ;
        RECT 217.230 185.520 217.490 185.840 ;
        RECT 216.770 184.500 217.030 184.820 ;
        RECT 215.850 183.820 216.110 184.140 ;
        RECT 215.910 179.040 216.050 183.820 ;
        RECT 217.290 181.420 217.430 185.520 ;
        RECT 217.690 183.480 217.950 183.800 ;
        RECT 217.230 181.100 217.490 181.420 ;
        RECT 216.300 180.565 216.580 180.935 ;
        RECT 216.310 180.420 216.570 180.565 ;
        RECT 217.230 180.420 217.490 180.740 ;
        RECT 217.290 180.255 217.430 180.420 ;
        RECT 217.220 179.885 217.500 180.255 ;
        RECT 217.750 179.575 217.890 183.480 ;
        RECT 217.680 179.205 217.960 179.575 ;
        RECT 215.850 178.720 216.110 179.040 ;
        RECT 218.210 178.780 218.350 186.880 ;
        RECT 218.610 186.540 218.870 186.860 ;
        RECT 217.290 178.640 218.350 178.780 ;
        RECT 214.530 177.960 215.590 178.100 ;
        RECT 215.850 178.040 216.110 178.360 ;
        RECT 214.530 176.290 214.670 177.960 ;
        RECT 215.380 177.165 215.660 177.535 ;
        RECT 215.450 176.290 215.590 177.165 ;
        RECT 215.910 176.660 216.050 178.040 ;
        RECT 215.850 176.340 216.110 176.660 ;
        RECT 216.370 176.430 216.970 176.570 ;
        RECT 216.370 176.290 216.510 176.430 ;
        RECT 208.940 130.365 209.220 176.290 ;
        RECT 209.860 130.945 210.140 176.290 ;
        RECT 210.780 131.525 211.060 176.290 ;
        RECT 211.700 132.105 211.980 176.290 ;
        RECT 212.620 132.685 212.900 176.290 ;
        RECT 213.540 133.265 213.820 176.290 ;
        RECT 214.460 133.845 214.740 176.290 ;
        RECT 215.380 134.425 215.660 176.290 ;
        RECT 216.300 135.005 216.580 176.290 ;
        RECT 216.830 175.300 216.970 176.430 ;
        RECT 217.290 176.290 217.430 178.640 ;
        RECT 217.690 178.040 217.950 178.360 ;
        RECT 217.750 176.320 217.890 178.040 ;
        RECT 218.670 177.535 218.810 186.540 ;
        RECT 219.530 185.520 219.790 185.840 ;
        RECT 219.070 184.160 219.330 184.480 ;
        RECT 219.130 179.575 219.270 184.160 ;
        RECT 219.060 179.205 219.340 179.575 ;
        RECT 219.590 178.360 219.730 185.520 ;
        RECT 219.530 178.040 219.790 178.360 ;
        RECT 218.600 177.165 218.880 177.535 ;
        RECT 218.210 176.430 218.810 176.570 ;
        RECT 216.770 174.980 217.030 175.300 ;
        RECT 217.220 135.585 217.500 176.290 ;
        RECT 217.690 176.000 217.950 176.320 ;
        RECT 218.210 176.290 218.350 176.430 ;
        RECT 218.140 136.165 218.420 176.290 ;
        RECT 218.670 175.640 218.810 176.430 ;
        RECT 219.130 176.430 219.730 176.570 ;
        RECT 219.130 176.290 219.270 176.430 ;
        RECT 218.610 175.320 218.870 175.640 ;
        RECT 219.060 136.745 219.340 176.290 ;
        RECT 219.590 175.980 219.730 176.430 ;
        RECT 220.050 176.290 220.190 186.880 ;
        RECT 220.450 185.860 220.710 186.180 ;
        RECT 220.510 177.680 220.650 185.860 ;
        RECT 222.290 185.520 222.550 185.840 ;
        RECT 221.370 184.160 221.630 184.480 ;
        RECT 221.430 178.700 221.570 184.160 ;
        RECT 222.350 181.420 222.490 185.520 ;
        RECT 224.650 184.140 224.790 189.520 ;
        RECT 230.570 189.260 230.830 189.580 ;
        RECT 225.050 188.920 225.310 189.240 ;
        RECT 228.270 188.920 228.530 189.240 ;
        RECT 229.190 188.920 229.450 189.240 ;
        RECT 225.110 187.540 225.250 188.920 ;
        RECT 227.350 188.240 227.610 188.560 ;
        RECT 225.050 187.220 225.310 187.540 ;
        RECT 227.410 186.520 227.550 188.240 ;
        RECT 227.810 186.540 228.070 186.860 ;
        RECT 227.350 186.200 227.610 186.520 ;
        RECT 225.510 185.860 225.770 186.180 ;
        RECT 224.590 183.820 224.850 184.140 ;
        RECT 223.660 183.285 223.940 183.655 ;
        RECT 224.580 183.285 224.860 183.655 ;
        RECT 222.750 181.780 223.010 182.100 ;
        RECT 222.290 181.100 222.550 181.420 ;
        RECT 221.830 180.760 222.090 181.080 ;
        RECT 221.890 180.255 222.030 180.760 ;
        RECT 221.820 179.885 222.100 180.255 ;
        RECT 221.370 178.380 221.630 178.700 ;
        RECT 220.450 177.360 220.710 177.680 ;
        RECT 220.910 177.360 221.170 177.680 ;
        RECT 220.970 176.290 221.110 177.360 ;
        RECT 221.430 176.320 221.570 178.380 ;
        RECT 221.890 176.600 222.490 176.740 ;
        RECT 219.530 175.660 219.790 175.980 ;
        RECT 219.980 137.325 220.260 176.290 ;
        RECT 220.900 137.905 221.180 176.290 ;
        RECT 221.370 176.000 221.630 176.320 ;
        RECT 221.890 176.290 222.030 176.600 ;
        RECT 222.350 176.320 222.490 176.600 ;
        RECT 221.820 138.485 222.100 176.290 ;
        RECT 222.290 176.000 222.550 176.320 ;
        RECT 222.810 176.290 222.950 181.780 ;
        RECT 223.210 180.760 223.470 181.080 ;
        RECT 223.270 178.215 223.410 180.760 ;
        RECT 223.200 177.845 223.480 178.215 ;
        RECT 223.730 176.290 223.870 183.285 ;
        RECT 224.650 183.120 224.790 183.285 ;
        RECT 224.130 182.800 224.390 183.120 ;
        RECT 224.590 182.800 224.850 183.120 ;
        RECT 224.190 181.080 224.330 182.800 ;
        RECT 224.130 180.760 224.390 181.080 ;
        RECT 225.570 180.740 225.710 185.860 ;
        RECT 225.970 183.480 226.230 183.800 ;
        RECT 225.510 180.420 225.770 180.740 ;
        RECT 226.030 178.360 226.170 183.480 ;
        RECT 227.340 183.285 227.620 183.655 ;
        RECT 226.430 180.080 226.690 180.400 ;
        RECT 226.490 178.895 226.630 180.080 ;
        RECT 226.420 178.525 226.700 178.895 ;
        RECT 224.590 178.100 224.850 178.360 ;
        RECT 225.970 178.215 226.230 178.360 ;
        RECT 224.590 178.040 225.710 178.100 ;
        RECT 224.650 177.960 225.710 178.040 ;
        RECT 225.570 177.590 225.710 177.960 ;
        RECT 225.960 177.845 226.240 178.215 ;
        RECT 227.410 177.590 227.550 183.285 ;
        RECT 227.870 181.615 228.010 186.540 ;
        RECT 227.800 181.245 228.080 181.615 ;
        RECT 227.810 180.935 228.070 181.080 ;
        RECT 227.800 180.565 228.080 180.935 ;
        RECT 227.810 180.080 228.070 180.400 ;
        RECT 225.570 177.450 226.170 177.590 ;
        RECT 224.650 176.430 225.250 176.570 ;
        RECT 225.500 176.485 225.780 176.855 ;
        RECT 226.030 176.660 226.170 177.450 ;
        RECT 226.490 177.450 227.550 177.590 ;
        RECT 227.870 177.535 228.010 180.080 ;
        RECT 228.330 179.380 228.470 188.920 ;
        RECT 229.250 188.160 229.390 188.920 ;
        RECT 229.650 188.580 229.910 188.900 ;
        RECT 228.790 188.020 229.390 188.160 ;
        RECT 228.270 179.060 228.530 179.380 ;
        RECT 228.790 178.780 228.930 188.020 ;
        RECT 229.190 185.520 229.450 185.840 ;
        RECT 229.250 184.820 229.390 185.520 ;
        RECT 229.190 184.500 229.450 184.820 ;
        RECT 229.190 183.480 229.450 183.800 ;
        RECT 229.250 182.100 229.390 183.480 ;
        RECT 229.190 181.780 229.450 182.100 ;
        RECT 229.710 179.460 229.850 188.580 ;
        RECT 230.630 187.735 230.770 189.260 ;
        RECT 231.030 188.580 231.290 188.900 ;
        RECT 230.560 187.365 230.840 187.735 ;
        RECT 230.110 184.500 230.370 184.820 ;
        RECT 230.170 183.655 230.310 184.500 ;
        RECT 230.570 184.160 230.830 184.480 ;
        RECT 230.100 183.285 230.380 183.655 ;
        RECT 230.110 182.800 230.370 183.120 ;
        RECT 228.330 178.640 228.930 178.780 ;
        RECT 229.250 179.320 229.850 179.460 ;
        RECT 224.650 176.290 224.790 176.430 ;
        RECT 222.740 139.065 223.020 176.290 ;
        RECT 223.660 139.645 223.940 176.290 ;
        RECT 224.580 140.225 224.860 176.290 ;
        RECT 225.110 176.175 225.250 176.430 ;
        RECT 225.570 176.290 225.710 176.485 ;
        RECT 225.970 176.340 226.230 176.660 ;
        RECT 226.490 176.290 226.630 177.450 ;
        RECT 227.800 177.165 228.080 177.535 ;
        RECT 227.340 176.485 227.620 176.855 ;
        RECT 227.410 176.290 227.550 176.485 ;
        RECT 228.330 176.290 228.470 178.640 ;
        RECT 229.250 176.290 229.390 179.320 ;
        RECT 230.170 178.700 230.310 182.800 ;
        RECT 230.630 179.380 230.770 184.160 ;
        RECT 230.570 179.060 230.830 179.380 ;
        RECT 230.110 178.380 230.370 178.700 ;
        RECT 229.650 178.040 229.910 178.360 ;
        RECT 225.040 175.805 225.320 176.175 ;
        RECT 225.500 140.805 225.780 176.290 ;
        RECT 226.420 141.385 226.700 176.290 ;
        RECT 227.340 141.965 227.620 176.290 ;
        RECT 228.260 142.545 228.540 176.290 ;
        RECT 229.180 143.125 229.460 176.290 ;
        RECT 229.710 175.300 229.850 178.040 ;
        RECT 230.100 177.845 230.380 178.215 ;
        RECT 230.170 176.290 230.310 177.845 ;
        RECT 231.090 176.290 231.230 188.580 ;
        RECT 231.550 181.340 231.690 189.600 ;
        RECT 232.470 187.540 232.610 190.960 ;
        RECT 232.410 187.220 232.670 187.540 ;
        RECT 232.860 187.365 233.140 187.735 ;
        RECT 236.150 187.540 236.290 199.800 ;
        RECT 232.930 186.860 233.070 187.365 ;
        RECT 236.090 187.220 236.350 187.540 ;
        RECT 232.870 186.540 233.130 186.860 ;
        RECT 233.780 186.685 234.060 187.055 ;
        RECT 233.790 186.540 234.050 186.685 ;
        RECT 236.090 186.540 236.350 186.860 ;
        RECT 231.950 185.860 232.210 186.180 ;
        RECT 232.010 181.500 232.150 185.860 ;
        RECT 235.170 185.520 235.430 185.840 ;
        RECT 234.240 184.645 234.520 185.015 ;
        RECT 234.250 184.500 234.510 184.645 ;
        RECT 234.250 183.480 234.510 183.800 ;
        RECT 233.330 183.140 233.590 183.460 ;
        RECT 232.400 182.605 232.680 182.975 ;
        RECT 232.870 182.800 233.130 183.120 ;
        RECT 232.470 182.100 232.610 182.605 ;
        RECT 232.930 182.295 233.070 182.800 ;
        RECT 232.410 181.780 232.670 182.100 ;
        RECT 232.860 181.925 233.140 182.295 ;
        RECT 232.010 181.420 233.070 181.500 ;
        RECT 232.010 181.360 233.130 181.420 ;
        RECT 231.490 181.020 231.750 181.340 ;
        RECT 232.870 181.100 233.130 181.360 ;
        RECT 232.410 180.760 232.670 181.080 ;
        RECT 231.480 179.205 231.760 179.575 ;
        RECT 232.470 179.380 232.610 180.760 ;
        RECT 231.490 179.060 231.750 179.205 ;
        RECT 232.410 179.060 232.670 179.380 ;
        RECT 232.930 178.895 233.070 181.100 ;
        RECT 232.860 178.525 233.140 178.895 ;
        RECT 232.410 178.040 232.670 178.360 ;
        RECT 229.650 174.980 229.910 175.300 ;
        RECT 230.100 143.705 230.380 176.290 ;
        RECT 231.020 144.285 231.300 176.290 ;
        RECT 232.470 175.640 232.610 178.040 ;
        RECT 233.390 176.855 233.530 183.140 ;
        RECT 233.790 178.040 234.050 178.360 ;
        RECT 233.320 176.485 233.600 176.855 ;
        RECT 233.850 175.980 233.990 178.040 ;
        RECT 234.310 176.175 234.450 183.480 ;
        RECT 234.700 181.245 234.980 181.615 ;
        RECT 234.770 179.380 234.910 181.245 ;
        RECT 234.710 179.060 234.970 179.380 ;
        RECT 235.230 176.660 235.370 185.520 ;
        RECT 235.630 182.800 235.890 183.120 ;
        RECT 235.690 180.255 235.830 182.800 ;
        RECT 235.620 179.885 235.900 180.255 ;
        RECT 236.150 178.215 236.290 186.540 ;
        RECT 236.540 186.005 236.820 186.375 ;
        RECT 236.610 181.080 236.750 186.005 ;
        RECT 236.550 180.760 236.810 181.080 ;
        RECT 236.080 177.845 236.360 178.215 ;
        RECT 236.550 178.040 236.810 178.360 ;
        RECT 235.170 176.340 235.430 176.660 ;
        RECT 236.610 176.320 236.750 178.040 ;
        RECT 233.790 175.660 234.050 175.980 ;
        RECT 234.240 175.805 234.520 176.175 ;
        RECT 236.550 176.000 236.810 176.320 ;
        RECT 232.410 175.320 232.670 175.640 ;
        RECT 231.020 144.005 309.205 144.285 ;
        RECT 230.100 143.425 306.905 143.705 ;
        RECT 229.180 142.845 304.605 143.125 ;
        RECT 228.260 142.265 302.305 142.545 ;
        RECT 227.340 141.685 300.005 141.965 ;
        RECT 226.420 141.105 297.705 141.385 ;
        RECT 225.500 140.525 295.405 140.805 ;
        RECT 224.580 139.945 293.105 140.225 ;
        RECT 223.660 139.365 290.805 139.645 ;
        RECT 222.740 138.785 288.505 139.065 ;
        RECT 221.820 138.205 286.205 138.485 ;
        RECT 220.900 137.625 283.905 137.905 ;
        RECT 219.980 137.045 281.605 137.325 ;
        RECT 219.060 136.465 279.305 136.745 ;
        RECT 218.140 135.885 277.005 136.165 ;
        RECT 217.220 135.305 274.705 135.585 ;
        RECT 216.300 134.725 272.405 135.005 ;
        RECT 215.380 134.145 270.105 134.425 ;
        RECT 214.460 133.565 267.805 133.845 ;
        RECT 213.540 132.985 265.505 133.265 ;
        RECT 212.620 132.405 263.205 132.685 ;
        RECT 211.700 131.825 260.905 132.105 ;
        RECT 210.780 131.245 258.605 131.525 ;
        RECT 209.860 130.665 256.305 130.945 ;
        RECT 208.940 130.085 254.005 130.365 ;
        RECT 208.020 129.505 251.705 129.785 ;
        RECT 207.100 128.925 249.405 129.205 ;
        RECT 206.180 128.345 247.105 128.625 ;
        RECT 205.260 127.765 244.805 128.045 ;
        RECT 204.340 127.185 242.505 127.465 ;
        RECT 203.420 126.605 240.205 126.885 ;
        RECT 202.500 126.025 237.905 126.305 ;
        RECT 201.580 125.445 235.605 125.725 ;
        RECT 200.660 124.865 233.305 125.145 ;
        RECT 199.740 124.285 231.005 124.565 ;
        RECT 198.820 123.705 228.705 123.985 ;
        RECT 197.900 123.125 226.405 123.405 ;
        RECT 196.980 122.545 224.105 122.825 ;
        RECT 196.060 121.965 221.805 122.245 ;
        RECT 195.140 121.385 219.505 121.665 ;
        RECT 194.220 120.805 217.205 121.085 ;
        RECT 193.300 120.225 214.905 120.505 ;
        RECT 192.380 119.645 212.605 119.925 ;
        RECT 191.460 119.065 210.305 119.345 ;
        RECT 190.540 118.485 208.005 118.765 ;
        RECT 189.620 117.905 205.705 118.185 ;
        RECT 188.700 117.325 203.405 117.605 ;
        RECT 187.780 116.745 201.105 117.025 ;
        RECT 186.860 116.165 198.805 116.445 ;
        RECT 185.940 115.585 196.505 115.865 ;
        RECT 185.020 115.005 194.205 115.285 ;
        RECT 184.100 114.425 191.905 114.705 ;
        RECT 183.180 113.845 189.605 114.125 ;
        RECT 182.260 113.265 187.305 113.545 ;
        RECT 181.340 112.685 185.005 112.965 ;
        RECT 180.420 112.105 182.705 112.385 ;
        RECT 179.500 111.525 180.405 111.805 ;
        RECT 177.825 109.225 178.105 111.525 ;
        RECT 180.125 109.225 180.405 111.525 ;
        RECT 182.425 109.225 182.705 112.105 ;
        RECT 184.725 109.225 185.005 112.685 ;
        RECT 187.025 109.225 187.305 113.265 ;
        RECT 189.325 109.225 189.605 113.845 ;
        RECT 191.625 109.225 191.905 114.425 ;
        RECT 193.925 109.225 194.205 115.005 ;
        RECT 196.225 109.225 196.505 115.585 ;
        RECT 198.525 109.225 198.805 116.165 ;
        RECT 200.825 109.225 201.105 116.745 ;
        RECT 203.125 109.225 203.405 117.325 ;
        RECT 205.425 109.225 205.705 117.905 ;
        RECT 207.725 109.225 208.005 118.485 ;
        RECT 210.025 109.225 210.305 119.065 ;
        RECT 212.325 109.225 212.605 119.645 ;
        RECT 214.625 109.225 214.905 120.225 ;
        RECT 216.925 109.225 217.205 120.805 ;
        RECT 219.225 109.225 219.505 121.385 ;
        RECT 221.525 109.225 221.805 121.965 ;
        RECT 223.825 109.225 224.105 122.545 ;
        RECT 226.125 109.225 226.405 123.125 ;
        RECT 228.425 109.225 228.705 123.705 ;
        RECT 230.725 109.225 231.005 124.285 ;
        RECT 233.025 109.225 233.305 124.865 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 164.095 100.635 164.235 109.225 ;
        RECT 164.495 105.075 164.755 105.395 ;
        RECT 164.035 100.315 164.295 100.635 ;
        RECT 164.035 93.350 164.295 93.495 ;
        RECT 164.025 92.980 164.305 93.350 ;
        RECT 146.290 88.455 148.395 92.555 ;
        RECT 146.290 83.775 148.395 87.875 ;
        RECT 146.290 77.925 148.395 83.195 ;
        RECT 146.290 73.245 148.395 77.345 ;
        RECT 146.290 68.565 148.395 72.665 ;
        RECT 164.555 70.375 164.695 105.075 ;
        RECT 166.395 103.355 166.535 109.225 ;
        RECT 168.175 106.775 168.435 107.095 ;
        RECT 166.795 105.075 167.055 105.395 ;
        RECT 166.335 103.035 166.595 103.355 ;
        RECT 165.875 102.015 166.135 102.335 ;
        RECT 165.415 96.575 165.675 96.895 ;
        RECT 164.955 94.195 165.215 94.515 ;
        RECT 165.015 70.715 165.155 94.195 ;
        RECT 165.475 92.135 165.615 96.575 ;
        RECT 165.415 91.815 165.675 92.135 ;
        RECT 165.475 88.735 165.615 91.815 ;
        RECT 165.935 89.755 166.075 102.015 ;
        RECT 166.335 99.635 166.595 99.955 ;
        RECT 165.875 89.435 166.135 89.755 ;
        RECT 165.415 88.415 165.675 88.735 ;
        RECT 165.935 86.355 166.075 89.435 ;
        RECT 165.875 86.035 166.135 86.355 ;
        RECT 165.935 78.195 166.075 86.035 ;
        RECT 166.395 84.315 166.535 99.635 ;
        RECT 166.335 83.995 166.595 84.315 ;
        RECT 165.875 77.875 166.135 78.195 ;
        RECT 164.955 70.395 165.215 70.715 ;
        RECT 164.495 70.055 164.755 70.375 ;
        RECT 146.290 63.885 148.395 67.985 ;
        RECT 164.555 65.275 164.695 70.055 ;
        RECT 166.855 70.035 166.995 105.075 ;
        RECT 168.235 104.715 168.375 106.775 ;
        RECT 168.175 104.395 168.435 104.715 ;
        RECT 168.695 102.755 168.835 109.225 ;
        RECT 169.095 105.075 169.355 105.395 ;
        RECT 168.235 102.615 168.835 102.755 ;
        RECT 167.255 99.295 167.515 99.615 ;
        RECT 167.315 94.515 167.455 99.295 ;
        RECT 168.235 97.915 168.375 102.615 ;
        RECT 168.635 101.675 168.895 101.995 ;
        RECT 168.695 97.915 168.835 101.675 ;
        RECT 168.175 97.595 168.435 97.915 ;
        RECT 168.635 97.595 168.895 97.915 ;
        RECT 167.255 94.425 167.515 94.515 ;
        RECT 167.255 94.285 167.915 94.425 ;
        RECT 167.255 94.195 167.515 94.285 ;
        RECT 167.255 90.455 167.515 90.775 ;
        RECT 167.315 86.355 167.455 90.455 ;
        RECT 167.775 86.355 167.915 94.285 ;
        RECT 167.255 86.035 167.515 86.355 ;
        RECT 167.715 86.035 167.975 86.355 ;
        RECT 167.775 83.975 167.915 86.035 ;
        RECT 167.715 83.655 167.975 83.975 ;
        RECT 166.795 69.715 167.055 70.035 ;
        RECT 168.635 68.695 168.895 69.015 ;
        RECT 168.695 67.655 168.835 68.695 ;
        RECT 168.635 67.335 168.895 67.655 ;
        RECT 164.495 64.955 164.755 65.275 ;
        RECT 169.155 63.575 169.295 105.075 ;
        RECT 170.015 102.355 170.275 102.675 ;
        RECT 170.075 101.995 170.215 102.355 ;
        RECT 170.015 101.675 170.275 101.995 ;
        RECT 170.075 100.295 170.215 101.675 ;
        RECT 170.015 99.975 170.275 100.295 ;
        RECT 170.075 94.855 170.215 99.975 ;
        RECT 170.995 97.995 171.135 109.225 ;
        RECT 171.855 107.455 172.115 107.775 ;
        RECT 171.915 104.375 172.055 107.455 ;
        RECT 172.315 107.115 172.575 107.435 ;
        RECT 172.375 105.395 172.515 107.115 ;
        RECT 173.295 106.075 173.435 109.225 ;
        RECT 173.235 105.755 173.495 106.075 ;
        RECT 173.695 105.475 173.955 105.735 ;
        RECT 172.835 105.415 173.955 105.475 ;
        RECT 172.835 105.395 173.895 105.415 ;
        RECT 172.315 105.075 172.575 105.395 ;
        RECT 172.775 105.335 173.895 105.395 ;
        RECT 172.775 105.075 173.035 105.335 ;
        RECT 174.615 105.075 174.875 105.395 ;
        RECT 175.075 105.075 175.335 105.395 ;
        RECT 171.855 104.055 172.115 104.375 ;
        RECT 174.675 101.655 174.815 105.075 ;
        RECT 174.155 101.335 174.415 101.655 ;
        RECT 174.615 101.335 174.875 101.655 ;
        RECT 170.535 97.855 171.135 97.995 ;
        RECT 170.535 97.575 170.675 97.855 ;
        RECT 170.475 97.255 170.735 97.575 ;
        RECT 170.015 94.535 170.275 94.855 ;
        RECT 172.315 94.535 172.575 94.855 ;
        RECT 172.375 94.095 172.515 94.535 ;
        RECT 171.915 93.955 172.515 94.095 ;
        RECT 171.915 89.415 172.055 93.955 ;
        RECT 172.315 91.475 172.575 91.795 ;
        RECT 171.855 89.095 172.115 89.415 ;
        RECT 171.915 85.335 172.055 89.095 ;
        RECT 172.375 88.735 172.515 91.475 ;
        RECT 172.315 88.415 172.575 88.735 ;
        RECT 171.855 85.015 172.115 85.335 ;
        RECT 170.935 82.975 171.195 83.295 ;
        RECT 170.995 81.595 171.135 82.975 ;
        RECT 170.935 81.275 171.195 81.595 ;
        RECT 172.375 80.915 172.515 88.415 ;
        RECT 174.215 88.055 174.355 101.335 ;
        RECT 175.135 100.715 175.275 105.075 ;
        RECT 175.595 105.055 175.735 109.225 ;
        RECT 177.895 107.095 178.035 109.225 ;
        RECT 177.835 106.775 178.095 107.095 ;
        RECT 176.915 105.075 177.175 105.395 ;
        RECT 175.535 104.735 175.795 105.055 ;
        RECT 175.535 104.055 175.795 104.375 ;
        RECT 175.595 103.355 175.735 104.055 ;
        RECT 175.535 103.035 175.795 103.355 ;
        RECT 176.975 102.755 177.115 105.075 ;
        RECT 179.675 104.735 179.935 105.055 ;
        RECT 177.645 103.520 179.185 103.890 ;
        RECT 177.375 103.035 177.635 103.355 ;
        RECT 177.435 102.755 177.575 103.035 ;
        RECT 176.975 102.615 177.575 102.755 ;
        RECT 176.915 101.335 177.175 101.655 ;
        RECT 174.675 100.575 175.275 100.715 ;
        RECT 174.675 91.455 174.815 100.575 ;
        RECT 176.975 97.430 177.115 101.335 ;
        RECT 179.735 99.615 179.875 104.735 ;
        RECT 180.195 104.715 180.335 109.225 ;
        RECT 182.495 107.345 182.635 109.225 ;
        RECT 184.795 107.775 184.935 109.225 ;
        RECT 184.735 107.455 184.995 107.775 ;
        RECT 182.495 107.205 183.095 107.345 ;
        RECT 180.945 106.240 182.485 106.610 ;
        RECT 180.595 105.075 180.855 105.395 ;
        RECT 180.135 104.395 180.395 104.715 ;
        RECT 179.675 99.295 179.935 99.615 ;
        RECT 177.645 98.080 179.185 98.450 ;
        RECT 176.905 97.060 177.185 97.430 ;
        RECT 179.735 97.235 179.875 99.295 ;
        RECT 176.455 96.575 176.715 96.895 ;
        RECT 175.075 95.895 175.335 96.215 ;
        RECT 175.535 95.895 175.795 96.215 ;
        RECT 175.135 93.235 175.275 95.895 ;
        RECT 175.595 94.175 175.735 95.895 ;
        RECT 175.535 93.855 175.795 94.175 ;
        RECT 175.135 93.095 176.195 93.235 ;
        RECT 174.615 91.135 174.875 91.455 ;
        RECT 176.055 90.775 176.195 93.095 ;
        RECT 176.515 91.705 176.655 96.575 ;
        RECT 176.975 96.555 177.115 97.060 ;
        RECT 179.675 96.915 179.935 97.235 ;
        RECT 176.915 96.235 177.175 96.555 ;
        RECT 180.135 96.235 180.395 96.555 ;
        RECT 179.675 95.895 179.935 96.215 ;
        RECT 177.645 92.640 179.185 93.010 ;
        RECT 179.735 91.875 179.875 95.895 ;
        RECT 180.195 95.195 180.335 96.235 ;
        RECT 180.135 94.875 180.395 95.195 ;
        RECT 179.275 91.735 179.875 91.875 ;
        RECT 176.515 91.565 177.575 91.705 ;
        RECT 176.915 90.795 177.175 91.115 ;
        RECT 175.075 90.455 175.335 90.775 ;
        RECT 175.995 90.455 176.255 90.775 ;
        RECT 175.135 89.415 175.275 90.455 ;
        RECT 176.975 89.415 177.115 90.795 ;
        RECT 175.075 89.095 175.335 89.415 ;
        RECT 176.915 89.095 177.175 89.415 ;
        RECT 177.435 89.075 177.575 91.565 ;
        RECT 177.375 88.755 177.635 89.075 ;
        RECT 179.275 88.735 179.415 91.735 ;
        RECT 180.655 90.515 180.795 105.075 ;
        RECT 180.945 100.800 182.485 101.170 ;
        RECT 182.955 100.635 183.095 107.205 ;
        RECT 184.735 106.775 184.995 107.095 ;
        RECT 183.355 105.075 183.615 105.395 ;
        RECT 182.895 100.315 183.155 100.635 ;
        RECT 183.415 100.035 183.555 105.075 ;
        RECT 184.275 104.055 184.535 104.375 ;
        RECT 184.335 100.635 184.475 104.055 ;
        RECT 184.275 100.315 184.535 100.635 ;
        RECT 182.955 99.895 183.555 100.035 ;
        RECT 180.945 95.360 182.485 95.730 ;
        RECT 180.195 90.375 180.795 90.515 ;
        RECT 179.675 88.755 179.935 89.075 ;
        RECT 179.215 88.415 179.475 88.735 ;
        RECT 174.155 87.735 174.415 88.055 ;
        RECT 176.915 87.735 177.175 88.055 ;
        RECT 174.215 87.035 174.355 87.735 ;
        RECT 174.155 86.715 174.415 87.035 ;
        RECT 176.975 85.675 177.115 87.735 ;
        RECT 177.645 87.200 179.185 87.570 ;
        RECT 179.735 87.035 179.875 88.755 ;
        RECT 179.675 86.715 179.935 87.035 ;
        RECT 176.915 85.355 177.175 85.675 ;
        RECT 172.775 83.995 173.035 84.315 ;
        RECT 172.315 80.595 172.575 80.915 ;
        RECT 172.835 80.235 172.975 83.995 ;
        RECT 176.915 83.655 177.175 83.975 ;
        RECT 174.155 80.935 174.415 81.255 ;
        RECT 172.775 79.915 173.035 80.235 ;
        RECT 173.235 75.155 173.495 75.475 ;
        RECT 173.295 73.435 173.435 75.155 ;
        RECT 173.695 74.475 173.955 74.795 ;
        RECT 173.235 73.115 173.495 73.435 ;
        RECT 171.855 71.415 172.115 71.735 ;
        RECT 171.915 69.015 172.055 71.415 ;
        RECT 172.315 69.715 172.575 70.035 ;
        RECT 171.855 68.695 172.115 69.015 ;
        RECT 172.375 66.975 172.515 69.715 ;
        RECT 173.295 67.995 173.435 73.115 ;
        RECT 173.235 67.675 173.495 67.995 ;
        RECT 172.315 66.655 172.575 66.975 ;
        RECT 173.295 64.595 173.435 67.675 ;
        RECT 173.755 67.655 173.895 74.475 ;
        RECT 174.215 72.415 174.355 80.935 ;
        RECT 175.075 80.595 175.335 80.915 ;
        RECT 174.155 72.095 174.415 72.415 ;
        RECT 173.695 67.335 173.955 67.655 ;
        RECT 173.235 64.275 173.495 64.595 ;
        RECT 173.235 63.595 173.495 63.915 ;
        RECT 146.290 58.035 148.395 63.305 ;
        RECT 169.095 63.255 169.355 63.575 ;
        RECT 169.155 62.555 169.295 63.255 ;
        RECT 169.095 62.235 169.355 62.555 ;
        RECT 173.295 62.215 173.435 63.595 ;
        RECT 173.235 61.895 173.495 62.215 ;
        RECT 164.955 61.555 165.215 61.875 ;
        RECT 164.035 60.710 164.295 60.855 ;
        RECT 164.025 60.340 164.305 60.710 ;
        RECT 146.290 53.355 148.395 57.455 ;
        RECT 165.015 57.115 165.155 61.555 ;
        RECT 175.135 61.275 175.275 80.595 ;
        RECT 176.455 79.915 176.715 80.235 ;
        RECT 175.995 79.575 176.255 79.895 ;
        RECT 175.535 68.695 175.795 69.015 ;
        RECT 176.055 68.925 176.195 79.575 ;
        RECT 176.515 72.415 176.655 79.915 ;
        RECT 176.975 78.195 177.115 83.655 ;
        RECT 177.645 81.760 179.185 82.130 ;
        RECT 180.195 81.790 180.335 90.375 ;
        RECT 180.945 89.920 182.485 90.290 ;
        RECT 180.595 89.435 180.855 89.755 ;
        RECT 180.125 81.420 180.405 81.790 ;
        RECT 179.675 80.595 179.935 80.915 ;
        RECT 179.735 78.195 179.875 80.595 ;
        RECT 180.195 80.235 180.335 81.420 ;
        RECT 180.135 79.915 180.395 80.235 ;
        RECT 180.655 78.535 180.795 89.435 ;
        RECT 182.955 89.155 183.095 99.895 ;
        RECT 183.815 99.635 184.075 99.955 ;
        RECT 183.355 91.135 183.615 91.455 ;
        RECT 183.415 89.755 183.555 91.135 ;
        RECT 183.355 89.435 183.615 89.755 ;
        RECT 183.875 89.270 184.015 99.635 ;
        RECT 184.275 96.575 184.535 96.895 ;
        RECT 184.335 94.515 184.475 96.575 ;
        RECT 184.275 94.195 184.535 94.515 ;
        RECT 182.955 89.015 183.555 89.155 ;
        RECT 180.945 84.480 182.485 84.850 ;
        RECT 182.895 79.915 183.155 80.235 ;
        RECT 180.945 79.040 182.485 79.410 ;
        RECT 182.955 78.875 183.095 79.915 ;
        RECT 182.895 78.555 183.155 78.875 ;
        RECT 180.595 78.215 180.855 78.535 ;
        RECT 176.915 77.875 177.175 78.195 ;
        RECT 179.675 77.875 179.935 78.195 ;
        RECT 176.975 76.155 177.115 77.875 ;
        RECT 177.645 76.320 179.185 76.690 ;
        RECT 176.915 75.835 177.175 76.155 ;
        RECT 176.975 74.795 177.115 75.835 ;
        RECT 179.735 75.475 179.875 77.875 ;
        RECT 180.135 76.855 180.395 77.175 ;
        RECT 179.675 75.155 179.935 75.475 ;
        RECT 176.915 74.475 177.175 74.795 ;
        RECT 176.975 72.755 177.115 74.475 ;
        RECT 177.375 74.135 177.635 74.455 ;
        RECT 176.915 72.435 177.175 72.755 ;
        RECT 176.455 72.095 176.715 72.415 ;
        RECT 177.435 71.735 177.575 74.135 ;
        RECT 177.375 71.645 177.635 71.735 ;
        RECT 176.975 71.505 177.635 71.645 ;
        RECT 176.455 68.925 176.715 69.015 ;
        RECT 176.055 68.785 176.715 68.925 ;
        RECT 176.455 68.695 176.715 68.785 ;
        RECT 175.595 65.275 175.735 68.695 ;
        RECT 175.535 64.955 175.795 65.275 ;
        RECT 175.995 63.255 176.255 63.575 ;
        RECT 176.055 62.215 176.195 63.255 ;
        RECT 175.995 61.895 176.255 62.215 ;
        RECT 175.135 61.135 175.735 61.275 ;
        RECT 175.075 60.535 175.335 60.855 ;
        RECT 172.775 58.155 173.035 58.475 ;
        RECT 164.955 56.795 165.215 57.115 ;
        RECT 172.835 56.775 172.975 58.155 ;
        RECT 172.775 56.455 173.035 56.775 ;
        RECT 174.615 56.455 174.875 56.775 ;
        RECT 173.695 55.775 173.955 56.095 ;
        RECT 167.255 55.095 167.515 55.415 ;
        RECT 167.315 53.715 167.455 55.095 ;
        RECT 173.755 53.715 173.895 55.775 ;
        RECT 167.255 53.395 167.515 53.715 ;
        RECT 173.695 53.395 173.955 53.715 ;
        RECT 165.875 53.055 166.135 53.375 ;
        RECT 172.775 53.055 173.035 53.375 ;
        RECT 146.290 48.675 148.395 52.775 ;
        RECT 165.935 50.655 166.075 53.055 ;
        RECT 172.835 50.995 172.975 53.055 ;
        RECT 172.775 50.675 173.035 50.995 ;
        RECT 174.675 50.655 174.815 56.455 ;
        RECT 175.135 50.995 175.275 60.535 ;
        RECT 175.595 56.095 175.735 61.135 ;
        RECT 175.985 58.300 176.265 58.670 ;
        RECT 176.055 57.115 176.195 58.300 ;
        RECT 175.995 56.795 176.255 57.115 ;
        RECT 176.515 56.435 176.655 68.695 ;
        RECT 176.975 59.495 177.115 71.505 ;
        RECT 177.375 71.415 177.635 71.505 ;
        RECT 177.645 70.880 179.185 71.250 ;
        RECT 177.825 69.860 178.105 70.230 ;
        RECT 177.895 69.695 178.035 69.860 ;
        RECT 179.675 69.715 179.935 70.035 ;
        RECT 177.835 69.375 178.095 69.695 ;
        RECT 177.645 65.440 179.185 65.810 ;
        RECT 179.735 64.595 179.875 69.715 ;
        RECT 179.675 64.275 179.935 64.595 ;
        RECT 180.195 64.255 180.335 76.855 ;
        RECT 180.655 75.475 180.795 78.215 ;
        RECT 181.515 77.875 181.775 78.195 ;
        RECT 181.045 77.340 181.325 77.710 ;
        RECT 180.595 75.155 180.855 75.475 ;
        RECT 181.115 74.795 181.255 77.340 ;
        RECT 181.575 77.175 181.715 77.875 ;
        RECT 183.415 77.710 183.555 89.015 ;
        RECT 183.805 88.900 184.085 89.270 ;
        RECT 184.795 87.115 184.935 106.775 ;
        RECT 186.575 104.965 186.835 105.055 ;
        RECT 187.095 104.965 187.235 109.225 ;
        RECT 186.575 104.825 187.235 104.965 ;
        RECT 186.575 104.735 186.835 104.825 ;
        RECT 188.415 104.735 188.675 105.055 ;
        RECT 185.655 102.015 185.915 102.335 ;
        RECT 185.195 99.975 185.455 100.295 ;
        RECT 184.335 86.975 184.935 87.115 ;
        RECT 183.815 82.975 184.075 83.295 ;
        RECT 183.875 78.875 184.015 82.975 ;
        RECT 184.335 80.915 184.475 86.975 ;
        RECT 185.255 86.695 185.395 99.975 ;
        RECT 185.715 96.555 185.855 102.015 ;
        RECT 188.475 101.995 188.615 104.735 ;
        RECT 189.395 103.355 189.535 109.225 ;
        RECT 191.695 106.155 191.835 109.225 ;
        RECT 191.235 106.015 191.835 106.155 ;
        RECT 193.995 106.075 194.135 109.225 ;
        RECT 191.235 105.735 191.375 106.015 ;
        RECT 193.935 105.755 194.195 106.075 ;
        RECT 191.175 105.415 191.435 105.735 ;
        RECT 192.555 105.415 192.815 105.735 ;
        RECT 189.795 104.735 190.055 105.055 ;
        RECT 189.335 103.035 189.595 103.355 ;
        RECT 188.415 101.675 188.675 101.995 ;
        RECT 188.875 101.675 189.135 101.995 ;
        RECT 188.475 99.615 188.615 101.675 ;
        RECT 186.115 99.295 186.375 99.615 ;
        RECT 188.415 99.295 188.675 99.615 ;
        RECT 185.655 96.235 185.915 96.555 ;
        RECT 185.715 95.195 185.855 96.235 ;
        RECT 186.175 96.215 186.315 99.295 ;
        RECT 187.495 96.915 187.755 97.235 ;
        RECT 187.035 96.575 187.295 96.895 ;
        RECT 186.115 95.895 186.375 96.215 ;
        RECT 185.655 94.875 185.915 95.195 ;
        RECT 186.175 94.030 186.315 95.895 ;
        RECT 186.105 93.660 186.385 94.030 ;
        RECT 186.115 93.175 186.375 93.495 ;
        RECT 186.175 91.115 186.315 93.175 ;
        RECT 186.115 90.795 186.375 91.115 ;
        RECT 185.195 86.375 185.455 86.695 ;
        RECT 184.275 80.595 184.535 80.915 ;
        RECT 183.815 78.555 184.075 78.875 ;
        RECT 183.345 77.340 183.625 77.710 ;
        RECT 181.515 76.855 181.775 77.175 ;
        RECT 182.895 75.155 183.155 75.475 ;
        RECT 181.055 74.475 181.315 74.795 ;
        RECT 180.945 73.600 182.485 73.970 ;
        RECT 182.955 72.755 183.095 75.155 ;
        RECT 183.875 73.395 184.015 78.555 ;
        RECT 183.415 73.255 184.015 73.395 ;
        RECT 182.895 72.435 183.155 72.755 ;
        RECT 181.055 72.095 181.315 72.415 ;
        RECT 181.115 69.355 181.255 72.095 ;
        RECT 181.055 69.035 181.315 69.355 ;
        RECT 180.945 68.160 182.485 68.530 ;
        RECT 181.055 67.675 181.315 67.995 ;
        RECT 181.115 66.975 181.255 67.675 ;
        RECT 181.515 67.335 181.775 67.655 ;
        RECT 181.055 66.655 181.315 66.975 ;
        RECT 181.055 65.975 181.315 66.295 ;
        RECT 181.115 65.275 181.255 65.975 ;
        RECT 181.055 64.955 181.315 65.275 ;
        RECT 181.575 64.935 181.715 67.335 ;
        RECT 182.895 66.655 183.155 66.975 ;
        RECT 181.515 64.615 181.775 64.935 ;
        RECT 180.135 63.935 180.395 64.255 ;
        RECT 180.195 62.555 180.335 63.935 ;
        RECT 180.945 62.720 182.485 63.090 ;
        RECT 180.135 62.235 180.395 62.555 ;
        RECT 179.675 61.555 179.935 61.875 ;
        RECT 180.135 61.555 180.395 61.875 ;
        RECT 177.645 60.000 179.185 60.370 ;
        RECT 179.735 59.495 179.875 61.555 ;
        RECT 176.915 59.175 177.175 59.495 ;
        RECT 179.675 59.175 179.935 59.495 ;
        RECT 175.995 56.115 176.255 56.435 ;
        RECT 176.455 56.115 176.715 56.435 ;
        RECT 179.215 56.345 179.475 56.435 ;
        RECT 179.735 56.345 179.875 59.175 ;
        RECT 179.215 56.205 179.875 56.345 ;
        RECT 179.215 56.115 179.475 56.205 ;
        RECT 175.535 55.775 175.795 56.095 ;
        RECT 175.595 53.115 175.735 55.775 ;
        RECT 176.055 54.055 176.195 56.115 ;
        RECT 179.735 55.415 179.875 56.205 ;
        RECT 179.675 55.095 179.935 55.415 ;
        RECT 177.645 54.560 179.185 54.930 ;
        RECT 175.995 53.910 176.255 54.055 ;
        RECT 175.985 53.540 176.265 53.910 ;
        RECT 176.915 53.395 177.175 53.715 ;
        RECT 175.595 52.975 176.195 53.115 ;
        RECT 175.535 52.375 175.795 52.695 ;
        RECT 175.595 51.675 175.735 52.375 ;
        RECT 175.535 51.355 175.795 51.675 ;
        RECT 175.075 50.675 175.335 50.995 ;
        RECT 165.875 50.335 166.135 50.655 ;
        RECT 174.615 50.335 174.875 50.655 ;
        RECT 146.290 43.995 148.395 48.095 ;
        RECT 165.935 45.215 166.075 50.335 ;
        RECT 172.315 46.935 172.575 47.255 ;
        RECT 165.875 44.895 166.135 45.215 ;
        RECT 143.435 41.655 145.540 42.245 ;
        RECT 143.835 41.605 145.135 41.655 ;
        RECT 7.065 36.430 8.665 39.630 ;
        RECT 10.170 37.965 74.550 38.965 ;
        RECT 79.810 38.185 127.975 39.285 ;
        RECT 10.170 35.440 74.550 36.940 ;
        RECT 79.810 36.685 127.975 37.785 ;
        RECT 79.810 35.185 127.975 36.285 ;
        RECT 136.295 35.805 138.400 39.905 ;
        RECT 146.290 38.145 148.395 43.415 ;
        RECT 165.935 42.495 166.075 44.895 ;
        RECT 165.875 42.175 166.135 42.495 ;
        RECT 10.170 33.440 74.550 34.940 ;
        RECT 79.810 33.685 127.975 34.785 ;
        RECT 10.170 31.440 74.550 32.940 ;
        RECT 79.810 32.185 127.975 33.285 ;
        RECT 79.810 30.685 127.975 31.785 ;
        RECT 136.295 31.125 138.400 35.225 ;
        RECT 146.290 33.465 148.395 37.565 ;
        RECT 165.935 34.675 166.075 42.175 ;
        RECT 167.715 39.455 167.975 39.775 ;
        RECT 169.555 39.455 169.815 39.775 ;
        RECT 165.875 34.355 166.135 34.675 ;
        RECT 143.640 32.295 145.745 32.885 ;
        RECT 167.775 31.955 167.915 39.455 ;
        RECT 169.615 38.075 169.755 39.455 ;
        RECT 169.555 37.755 169.815 38.075 ;
        RECT 170.935 34.015 171.195 34.335 ;
        RECT 167.715 31.635 167.975 31.955 ;
        RECT 167.255 30.955 167.515 31.275 ;
        RECT 10.170 28.035 74.550 30.415 ;
        RECT 79.810 28.165 127.975 30.285 ;
        RECT 138.950 29.955 141.055 30.545 ;
        RECT 167.315 29.915 167.455 30.955 ;
        RECT 167.255 29.595 167.515 29.915 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 164.035 28.070 164.295 28.215 ;
        RECT 10.170 25.510 74.550 27.010 ;
        RECT 79.810 26.665 127.975 27.765 ;
        RECT 164.025 27.700 164.305 28.070 ;
        RECT 170.995 27.195 171.135 34.015 ;
        RECT 172.375 29.235 172.515 46.935 ;
        RECT 175.135 46.235 175.275 50.675 ;
        RECT 176.055 47.935 176.195 52.975 ;
        RECT 176.975 51.675 177.115 53.395 ;
        RECT 180.195 53.375 180.335 61.555 ;
        RECT 181.515 59.175 181.775 59.495 ;
        RECT 181.575 58.815 181.715 59.175 ;
        RECT 181.515 58.495 181.775 58.815 ;
        RECT 182.955 58.135 183.095 66.655 ;
        RECT 183.415 59.155 183.555 73.255 ;
        RECT 183.815 69.550 184.075 69.695 ;
        RECT 183.805 69.180 184.085 69.550 ;
        RECT 183.355 58.835 183.615 59.155 ;
        RECT 182.895 57.815 183.155 58.135 ;
        RECT 180.945 57.280 182.485 57.650 ;
        RECT 180.595 56.115 180.855 56.435 ;
        RECT 180.135 53.055 180.395 53.375 ;
        RECT 180.655 53.035 180.795 56.115 ;
        RECT 183.875 55.155 184.015 69.180 ;
        RECT 184.335 66.295 184.475 80.595 ;
        RECT 185.255 80.575 185.395 86.375 ;
        RECT 186.175 83.975 186.315 90.795 ;
        RECT 186.575 88.755 186.835 89.075 ;
        RECT 186.115 83.655 186.375 83.975 ;
        RECT 185.195 80.255 185.455 80.575 ;
        RECT 186.635 78.275 186.775 88.755 ;
        RECT 187.095 88.735 187.235 96.575 ;
        RECT 187.035 88.590 187.295 88.735 ;
        RECT 187.025 88.220 187.305 88.590 ;
        RECT 187.035 85.695 187.295 86.015 ;
        RECT 187.095 81.255 187.235 85.695 ;
        RECT 187.035 80.935 187.295 81.255 ;
        RECT 187.555 78.275 187.695 96.915 ;
        RECT 187.955 95.895 188.215 96.215 ;
        RECT 188.015 91.795 188.155 95.895 ;
        RECT 187.955 91.475 188.215 91.795 ;
        RECT 187.955 90.455 188.215 90.775 ;
        RECT 188.015 88.055 188.155 90.455 ;
        RECT 187.955 87.735 188.215 88.055 ;
        RECT 188.015 86.695 188.155 87.735 ;
        RECT 187.955 86.375 188.215 86.695 ;
        RECT 188.475 86.355 188.615 99.295 ;
        RECT 188.935 97.915 189.075 101.675 ;
        RECT 189.855 100.635 189.995 104.735 ;
        RECT 191.175 101.675 191.435 101.995 ;
        RECT 189.795 100.315 190.055 100.635 ;
        RECT 191.235 100.295 191.375 101.675 ;
        RECT 190.255 99.975 190.515 100.295 ;
        RECT 191.175 99.975 191.435 100.295 ;
        RECT 188.875 97.595 189.135 97.915 ;
        RECT 190.315 96.750 190.455 99.975 ;
        RECT 190.245 96.380 190.525 96.750 ;
        RECT 190.315 96.215 190.455 96.380 ;
        RECT 190.255 95.895 190.515 96.215 ;
        RECT 191.235 95.195 191.375 99.975 ;
        RECT 192.095 98.615 192.355 98.935 ;
        RECT 192.155 97.235 192.295 98.615 ;
        RECT 192.095 96.915 192.355 97.235 ;
        RECT 191.635 96.575 191.895 96.895 ;
        RECT 191.175 94.875 191.435 95.195 ;
        RECT 189.335 94.195 189.595 94.515 ;
        RECT 188.865 93.660 189.145 94.030 ;
        RECT 188.415 86.035 188.675 86.355 ;
        RECT 188.935 83.975 189.075 93.660 ;
        RECT 189.395 89.415 189.535 94.195 ;
        RECT 191.235 91.115 191.375 94.875 ;
        RECT 191.695 91.705 191.835 96.575 ;
        RECT 192.155 95.195 192.295 96.915 ;
        RECT 192.095 94.875 192.355 95.195 ;
        RECT 192.615 94.855 192.755 105.415 ;
        RECT 196.295 103.355 196.435 109.225 ;
        RECT 198.595 103.355 198.735 109.225 ;
        RECT 198.995 105.075 199.255 105.395 ;
        RECT 196.235 103.035 196.495 103.355 ;
        RECT 198.535 103.035 198.795 103.355 ;
        RECT 197.615 102.015 197.875 102.335 ;
        RECT 196.235 101.335 196.495 101.655 ;
        RECT 194.385 99.100 194.665 99.470 ;
        RECT 193.015 98.615 193.275 98.935 ;
        RECT 192.555 94.535 192.815 94.855 ;
        RECT 192.095 91.705 192.355 91.795 ;
        RECT 191.695 91.565 192.355 91.705 ;
        RECT 192.095 91.475 192.355 91.565 ;
        RECT 192.155 91.310 192.295 91.475 ;
        RECT 191.175 90.795 191.435 91.115 ;
        RECT 191.635 90.795 191.895 91.115 ;
        RECT 192.085 90.940 192.365 91.310 ;
        RECT 189.335 89.095 189.595 89.415 ;
        RECT 191.175 89.095 191.435 89.415 ;
        RECT 189.335 85.755 189.595 86.015 ;
        RECT 189.335 85.695 189.995 85.755 ;
        RECT 189.395 85.615 189.995 85.695 ;
        RECT 189.335 85.015 189.595 85.335 ;
        RECT 188.875 83.655 189.135 83.975 ;
        RECT 186.175 78.135 186.775 78.275 ;
        RECT 187.095 78.195 187.695 78.275 ;
        RECT 187.035 78.135 187.695 78.195 ;
        RECT 184.735 77.535 184.995 77.855 ;
        RECT 184.795 72.270 184.935 77.535 ;
        RECT 184.725 71.900 185.005 72.270 ;
        RECT 184.795 66.635 184.935 71.900 ;
        RECT 185.655 70.285 185.915 70.375 ;
        RECT 186.175 70.285 186.315 78.135 ;
        RECT 187.035 77.875 187.295 78.135 ;
        RECT 186.575 77.195 186.835 77.515 ;
        RECT 186.635 73.095 186.775 77.195 ;
        RECT 186.575 72.775 186.835 73.095 ;
        RECT 187.555 70.715 187.695 78.135 ;
        RECT 187.955 77.875 188.215 78.195 ;
        RECT 188.015 72.415 188.155 77.875 ;
        RECT 189.395 77.855 189.535 85.015 ;
        RECT 189.855 83.635 189.995 85.615 ;
        RECT 189.795 83.315 190.055 83.635 ;
        RECT 189.335 77.535 189.595 77.855 ;
        RECT 188.875 74.195 189.135 74.455 ;
        RECT 188.475 74.135 189.135 74.195 ;
        RECT 188.475 74.055 189.075 74.135 ;
        RECT 187.955 72.095 188.215 72.415 ;
        RECT 187.035 70.395 187.295 70.715 ;
        RECT 187.495 70.395 187.755 70.715 ;
        RECT 185.655 70.145 186.315 70.285 ;
        RECT 185.655 70.055 185.915 70.145 ;
        RECT 185.195 69.375 185.455 69.695 ;
        RECT 184.735 66.315 184.995 66.635 ;
        RECT 184.275 65.975 184.535 66.295 ;
        RECT 184.275 61.555 184.535 61.875 ;
        RECT 184.335 58.815 184.475 61.555 ;
        RECT 184.735 61.215 184.995 61.535 ;
        RECT 184.795 59.495 184.935 61.215 ;
        RECT 184.735 59.175 184.995 59.495 ;
        RECT 184.275 58.495 184.535 58.815 ;
        RECT 184.335 57.115 184.475 58.495 ;
        RECT 184.795 58.135 184.935 59.175 ;
        RECT 184.735 57.815 184.995 58.135 ;
        RECT 184.275 56.795 184.535 57.115 ;
        RECT 185.255 56.435 185.395 69.375 ;
        RECT 185.715 67.510 185.855 70.055 ;
        RECT 187.095 69.695 187.235 70.395 ;
        RECT 186.115 69.550 186.375 69.695 ;
        RECT 186.105 69.180 186.385 69.550 ;
        RECT 187.035 69.375 187.295 69.695 ;
        RECT 185.645 67.140 185.925 67.510 ;
        RECT 186.175 66.150 186.315 69.180 ;
        RECT 187.555 67.655 187.695 70.395 ;
        RECT 187.495 67.335 187.755 67.655 ;
        RECT 188.015 67.315 188.155 72.095 ;
        RECT 188.475 70.715 188.615 74.055 ;
        RECT 188.875 73.115 189.135 73.435 ;
        RECT 188.935 72.950 189.075 73.115 ;
        RECT 188.865 72.580 189.145 72.950 ;
        RECT 188.415 70.395 188.675 70.715 ;
        RECT 187.955 66.995 188.215 67.315 ;
        RECT 186.105 65.780 186.385 66.150 ;
        RECT 186.575 65.975 186.835 66.295 ;
        RECT 188.875 65.975 189.135 66.295 ;
        RECT 186.635 65.275 186.775 65.975 ;
        RECT 186.575 64.955 186.835 65.275 ;
        RECT 185.655 64.615 185.915 64.935 ;
        RECT 185.715 57.310 185.855 64.615 ;
        RECT 186.635 64.255 186.775 64.955 ;
        RECT 188.935 64.595 189.075 65.975 ;
        RECT 188.875 64.275 189.135 64.595 ;
        RECT 186.575 63.935 186.835 64.255 ;
        RECT 189.395 62.555 189.535 77.535 ;
        RECT 188.415 62.235 188.675 62.555 ;
        RECT 189.335 62.235 189.595 62.555 ;
        RECT 188.475 61.875 188.615 62.235 ;
        RECT 188.415 61.555 188.675 61.875 ;
        RECT 189.335 61.555 189.595 61.875 ;
        RECT 187.495 61.215 187.755 61.535 ;
        RECT 186.115 60.535 186.375 60.855 ;
        RECT 186.175 58.825 186.315 60.535 ;
        RECT 187.035 59.175 187.295 59.495 ;
        RECT 186.115 58.505 186.375 58.825 ;
        RECT 186.575 58.495 186.835 58.815 ;
        RECT 185.645 56.940 185.925 57.310 ;
        RECT 186.635 57.115 186.775 58.495 ;
        RECT 186.575 56.795 186.835 57.115 ;
        RECT 185.195 56.115 185.455 56.435 ;
        RECT 186.115 56.115 186.375 56.435 ;
        RECT 184.735 55.435 184.995 55.755 ;
        RECT 183.415 55.015 184.015 55.155 ;
        RECT 183.415 54.395 183.555 55.015 ;
        RECT 183.355 54.075 183.615 54.395 ;
        RECT 183.805 54.220 184.085 54.590 ;
        RECT 180.595 52.715 180.855 53.035 ;
        RECT 180.945 51.840 182.485 52.210 ;
        RECT 176.915 51.355 177.175 51.675 ;
        RECT 176.455 50.335 176.715 50.655 ;
        RECT 176.515 48.955 176.655 50.335 ;
        RECT 176.455 48.635 176.715 48.955 ;
        RECT 176.975 48.275 177.115 51.355 ;
        RECT 178.755 51.245 179.015 51.335 ;
        RECT 178.755 51.105 179.875 51.245 ;
        RECT 178.755 51.015 179.015 51.105 ;
        RECT 177.645 49.120 179.185 49.490 ;
        RECT 179.735 48.615 179.875 51.105 ;
        RECT 183.415 49.035 183.555 54.075 ;
        RECT 183.875 54.055 184.015 54.220 ;
        RECT 183.815 53.735 184.075 54.055 ;
        RECT 184.275 53.735 184.535 54.055 ;
        RECT 183.875 50.655 184.015 53.735 ;
        RECT 184.335 52.695 184.475 53.735 ;
        RECT 184.795 52.695 184.935 55.435 ;
        RECT 186.175 54.055 186.315 56.115 ;
        RECT 187.095 54.395 187.235 59.175 ;
        RECT 187.555 58.815 187.695 61.215 ;
        RECT 188.475 59.155 188.615 61.555 ;
        RECT 188.875 60.875 189.135 61.195 ;
        RECT 188.935 59.495 189.075 60.875 ;
        RECT 188.875 59.175 189.135 59.495 ;
        RECT 188.415 58.835 188.675 59.155 ;
        RECT 187.495 58.495 187.755 58.815 ;
        RECT 187.035 54.075 187.295 54.395 ;
        RECT 186.115 53.735 186.375 54.055 ;
        RECT 187.035 53.055 187.295 53.375 ;
        RECT 184.275 52.375 184.535 52.695 ;
        RECT 184.735 52.375 184.995 52.695 ;
        RECT 183.815 50.335 184.075 50.655 ;
        RECT 182.495 48.895 183.555 49.035 ;
        RECT 179.675 48.295 179.935 48.615 ;
        RECT 176.915 47.955 177.175 48.275 ;
        RECT 182.495 47.935 182.635 48.895 ;
        RECT 183.355 47.955 183.615 48.275 ;
        RECT 175.995 47.615 176.255 47.935 ;
        RECT 182.435 47.615 182.695 47.935 ;
        RECT 180.595 47.275 180.855 47.595 ;
        RECT 179.215 46.935 179.475 47.255 ;
        RECT 175.075 45.915 175.335 46.235 ;
        RECT 175.135 44.535 175.275 45.915 ;
        RECT 179.275 45.215 179.415 46.935 ;
        RECT 180.655 45.215 180.795 47.275 ;
        RECT 182.895 46.935 183.155 47.255 ;
        RECT 180.945 46.400 182.485 46.770 ;
        RECT 182.955 46.235 183.095 46.935 ;
        RECT 182.895 45.915 183.155 46.235 ;
        RECT 179.215 44.895 179.475 45.215 ;
        RECT 180.595 44.895 180.855 45.215 ;
        RECT 175.075 44.215 175.335 44.535 ;
        RECT 175.135 42.835 175.275 44.215 ;
        RECT 177.645 43.680 179.185 44.050 ;
        RECT 175.075 42.515 175.335 42.835 ;
        RECT 172.775 42.175 173.035 42.495 ;
        RECT 172.835 39.775 172.975 42.175 ;
        RECT 177.375 41.835 177.635 42.155 ;
        RECT 175.535 41.495 175.795 41.815 ;
        RECT 172.775 39.455 173.035 39.775 ;
        RECT 172.835 34.675 172.975 39.455 ;
        RECT 175.595 38.075 175.735 41.495 ;
        RECT 177.435 40.795 177.575 41.835 ;
        RECT 177.375 40.475 177.635 40.795 ;
        RECT 175.995 39.455 176.255 39.775 ;
        RECT 175.535 37.755 175.795 38.075 ;
        RECT 176.055 36.715 176.195 39.455 ;
        RECT 176.915 38.775 177.175 39.095 ;
        RECT 175.995 36.395 176.255 36.715 ;
        RECT 176.455 36.395 176.715 36.715 ;
        RECT 174.615 36.055 174.875 36.375 ;
        RECT 172.775 34.355 173.035 34.675 ;
        RECT 172.835 31.615 172.975 34.355 ;
        RECT 174.675 31.955 174.815 36.055 ;
        RECT 176.055 35.355 176.195 36.395 ;
        RECT 175.995 35.035 176.255 35.355 ;
        RECT 175.995 33.675 176.255 33.995 ;
        RECT 174.615 31.635 174.875 31.955 ;
        RECT 172.775 31.295 173.035 31.615 ;
        RECT 175.535 30.615 175.795 30.935 ;
        RECT 172.315 28.915 172.575 29.235 ;
        RECT 174.615 28.575 174.875 28.895 ;
        RECT 174.675 27.195 174.815 28.575 ;
        RECT 170.935 26.875 171.195 27.195 ;
        RECT 174.615 26.875 174.875 27.195 ;
        RECT 175.595 26.515 175.735 30.615 ;
        RECT 176.055 29.235 176.195 33.675 ;
        RECT 176.515 31.955 176.655 36.395 ;
        RECT 176.975 34.675 177.115 38.775 ;
        RECT 177.645 38.240 179.185 38.610 ;
        RECT 178.755 36.735 179.015 37.055 ;
        RECT 178.815 35.355 178.955 36.735 ;
        RECT 180.655 36.375 180.795 44.895 ;
        RECT 180.945 40.960 182.485 41.330 ;
        RECT 183.415 39.775 183.555 47.955 ;
        RECT 184.335 47.935 184.475 52.375 ;
        RECT 184.795 51.335 184.935 52.375 ;
        RECT 184.735 51.015 184.995 51.335 ;
        RECT 184.275 47.615 184.535 47.935 ;
        RECT 183.815 45.235 184.075 45.555 ;
        RECT 183.875 42.155 184.015 45.235 ;
        RECT 183.815 41.835 184.075 42.155 ;
        RECT 183.875 40.455 184.015 41.835 ;
        RECT 184.335 41.815 184.475 47.615 ;
        RECT 184.795 47.595 184.935 51.015 ;
        RECT 185.655 50.335 185.915 50.655 ;
        RECT 185.715 48.955 185.855 50.335 ;
        RECT 187.095 50.315 187.235 53.055 ;
        RECT 187.555 51.675 187.695 58.495 ;
        RECT 188.875 57.815 189.135 58.135 ;
        RECT 187.955 56.795 188.215 57.115 ;
        RECT 188.015 55.415 188.155 56.795 ;
        RECT 188.935 56.095 189.075 57.815 ;
        RECT 188.875 55.775 189.135 56.095 ;
        RECT 187.955 55.095 188.215 55.415 ;
        RECT 187.955 53.055 188.215 53.375 ;
        RECT 187.495 51.355 187.755 51.675 ;
        RECT 188.015 50.655 188.155 53.055 ;
        RECT 187.955 50.335 188.215 50.655 ;
        RECT 187.035 49.995 187.295 50.315 ;
        RECT 185.655 48.635 185.915 48.955 ;
        RECT 184.735 47.275 184.995 47.595 ;
        RECT 185.195 44.895 185.455 45.215 ;
        RECT 185.255 43.515 185.395 44.895 ;
        RECT 185.655 44.215 185.915 44.535 ;
        RECT 185.195 43.195 185.455 43.515 ;
        RECT 184.275 41.495 184.535 41.815 ;
        RECT 184.335 40.795 184.475 41.495 ;
        RECT 185.715 40.795 185.855 44.215 ;
        RECT 187.095 41.815 187.235 49.995 ;
        RECT 187.495 44.555 187.755 44.875 ;
        RECT 187.035 41.495 187.295 41.815 ;
        RECT 184.275 40.475 184.535 40.795 ;
        RECT 185.655 40.475 185.915 40.795 ;
        RECT 187.095 40.455 187.235 41.495 ;
        RECT 183.815 40.135 184.075 40.455 ;
        RECT 187.035 40.135 187.295 40.455 ;
        RECT 183.355 39.455 183.615 39.775 ;
        RECT 180.595 36.055 180.855 36.375 ;
        RECT 180.945 35.520 182.485 35.890 ;
        RECT 178.755 35.035 179.015 35.355 ;
        RECT 183.875 35.015 184.015 40.135 ;
        RECT 186.115 39.455 186.375 39.775 ;
        RECT 184.275 39.115 184.535 39.435 ;
        RECT 184.335 37.055 184.475 39.115 ;
        RECT 185.655 38.775 185.915 39.095 ;
        RECT 185.715 37.395 185.855 38.775 ;
        RECT 186.175 38.075 186.315 39.455 ;
        RECT 186.115 37.755 186.375 38.075 ;
        RECT 185.655 37.075 185.915 37.395 ;
        RECT 184.275 36.735 184.535 37.055 ;
        RECT 183.815 34.695 184.075 35.015 ;
        RECT 176.915 34.355 177.175 34.675 ;
        RECT 177.645 32.800 179.185 33.170 ;
        RECT 184.335 32.295 184.475 36.735 ;
        RECT 185.195 36.055 185.455 36.375 ;
        RECT 184.275 31.975 184.535 32.295 ;
        RECT 176.455 31.635 176.715 31.955 ;
        RECT 178.755 31.635 179.015 31.955 ;
        RECT 176.515 29.915 176.655 31.635 ;
        RECT 176.915 31.295 177.175 31.615 ;
        RECT 176.455 29.595 176.715 29.915 ;
        RECT 175.995 28.915 176.255 29.235 ;
        RECT 176.975 26.515 177.115 31.295 ;
        RECT 178.815 28.895 178.955 31.635 ;
        RECT 180.595 30.615 180.855 30.935 ;
        RECT 180.655 29.575 180.795 30.615 ;
        RECT 180.945 30.080 182.485 30.450 ;
        RECT 180.595 29.255 180.855 29.575 ;
        RECT 185.255 28.895 185.395 36.055 ;
        RECT 186.175 34.925 186.315 37.755 ;
        RECT 185.715 34.785 186.315 34.925 ;
        RECT 185.715 29.575 185.855 34.785 ;
        RECT 186.575 34.695 186.835 35.015 ;
        RECT 186.115 34.015 186.375 34.335 ;
        RECT 186.175 29.915 186.315 34.015 ;
        RECT 186.635 31.275 186.775 34.695 ;
        RECT 187.555 34.675 187.695 44.555 ;
        RECT 188.015 44.535 188.155 50.335 ;
        RECT 189.395 45.555 189.535 61.555 ;
        RECT 189.855 57.115 189.995 83.315 ;
        RECT 190.715 82.975 190.975 83.295 ;
        RECT 190.775 80.430 190.915 82.975 ;
        RECT 190.705 80.060 190.985 80.430 ;
        RECT 190.715 75.835 190.975 76.155 ;
        RECT 190.255 72.950 190.515 73.095 ;
        RECT 190.245 72.580 190.525 72.950 ;
        RECT 190.255 70.395 190.515 70.715 ;
        RECT 190.315 70.230 190.455 70.395 ;
        RECT 190.245 69.860 190.525 70.230 ;
        RECT 190.775 70.035 190.915 75.835 ;
        RECT 190.715 69.715 190.975 70.035 ;
        RECT 190.775 69.550 190.915 69.715 ;
        RECT 190.705 69.180 190.985 69.550 ;
        RECT 190.255 68.695 190.515 69.015 ;
        RECT 190.315 63.575 190.455 68.695 ;
        RECT 190.705 67.140 190.985 67.510 ;
        RECT 190.715 66.995 190.975 67.140 ;
        RECT 190.715 66.315 190.975 66.635 ;
        RECT 190.255 63.255 190.515 63.575 ;
        RECT 190.775 59.155 190.915 66.315 ;
        RECT 191.235 62.555 191.375 89.095 ;
        RECT 191.695 89.075 191.835 90.795 ;
        RECT 191.635 88.755 191.895 89.075 ;
        RECT 191.635 80.255 191.895 80.575 ;
        RECT 191.695 75.475 191.835 80.255 ;
        RECT 191.635 75.155 191.895 75.475 ;
        RECT 191.695 73.095 191.835 75.155 ;
        RECT 192.615 74.455 192.755 94.535 ;
        RECT 193.075 94.515 193.215 98.615 ;
        RECT 194.455 97.575 194.595 99.100 ;
        RECT 194.845 97.740 195.125 98.110 ;
        RECT 194.395 97.255 194.655 97.575 ;
        RECT 193.015 94.195 193.275 94.515 ;
        RECT 194.455 94.175 194.595 97.255 ;
        RECT 194.915 96.215 195.055 97.740 ;
        RECT 196.295 96.895 196.435 101.335 ;
        RECT 196.235 96.575 196.495 96.895 ;
        RECT 194.855 95.895 195.115 96.215 ;
        RECT 194.395 93.855 194.655 94.175 ;
        RECT 194.915 93.495 195.055 95.895 ;
        RECT 194.855 93.175 195.115 93.495 ;
        RECT 193.475 92.155 193.735 92.475 ;
        RECT 193.535 89.415 193.675 92.155 ;
        RECT 195.315 91.135 195.575 91.455 ;
        RECT 195.775 91.135 196.035 91.455 ;
        RECT 193.475 89.095 193.735 89.415 ;
        RECT 193.015 86.035 193.275 86.355 ;
        RECT 193.075 83.635 193.215 86.035 ;
        RECT 193.535 86.015 193.675 89.095 ;
        RECT 195.375 88.735 195.515 91.135 ;
        RECT 195.835 89.755 195.975 91.135 ;
        RECT 195.775 89.435 196.035 89.755 ;
        RECT 195.775 88.755 196.035 89.075 ;
        RECT 195.315 88.415 195.575 88.735 ;
        RECT 194.855 86.375 195.115 86.695 ;
        RECT 194.915 86.015 195.055 86.375 ;
        RECT 193.475 85.695 193.735 86.015 ;
        RECT 194.855 85.695 195.115 86.015 ;
        RECT 193.475 83.655 193.735 83.975 ;
        RECT 193.015 83.315 193.275 83.635 ;
        RECT 193.535 78.535 193.675 83.655 ;
        RECT 194.395 80.935 194.655 81.255 ;
        RECT 193.935 79.915 194.195 80.235 ;
        RECT 193.995 78.875 194.135 79.915 ;
        RECT 193.935 78.555 194.195 78.875 ;
        RECT 193.475 78.215 193.735 78.535 ;
        RECT 192.555 74.135 192.815 74.455 ;
        RECT 192.095 73.115 192.355 73.435 ;
        RECT 191.635 72.775 191.895 73.095 ;
        RECT 192.155 70.375 192.295 73.115 ;
        RECT 193.535 72.755 193.675 78.215 ;
        RECT 193.995 77.175 194.135 78.555 ;
        RECT 194.455 77.855 194.595 80.935 ;
        RECT 194.395 77.535 194.655 77.855 ;
        RECT 193.935 76.855 194.195 77.175 ;
        RECT 194.395 74.475 194.655 74.795 ;
        RECT 194.455 73.435 194.595 74.475 ;
        RECT 194.395 73.115 194.655 73.435 ;
        RECT 193.475 72.435 193.735 72.755 ;
        RECT 192.095 70.055 192.355 70.375 ;
        RECT 192.545 65.100 192.825 65.470 ;
        RECT 191.175 62.235 191.435 62.555 ;
        RECT 191.635 60.535 191.895 60.855 ;
        RECT 191.695 59.595 191.835 60.535 ;
        RECT 191.175 59.175 191.435 59.495 ;
        RECT 191.695 59.455 192.295 59.595 ;
        RECT 190.715 58.835 190.975 59.155 ;
        RECT 190.255 58.155 190.515 58.475 ;
        RECT 189.795 56.795 190.055 57.115 ;
        RECT 190.315 50.315 190.455 58.155 ;
        RECT 191.235 56.435 191.375 59.175 ;
        RECT 192.155 58.815 192.295 59.455 ;
        RECT 192.095 58.495 192.355 58.815 ;
        RECT 192.615 58.670 192.755 65.100 ;
        RECT 193.015 64.275 193.275 64.595 ;
        RECT 191.175 56.115 191.435 56.435 ;
        RECT 192.155 56.095 192.295 58.495 ;
        RECT 192.545 58.300 192.825 58.670 ;
        RECT 190.715 55.775 190.975 56.095 ;
        RECT 192.095 55.775 192.355 56.095 ;
        RECT 190.775 53.285 190.915 55.775 ;
        RECT 192.155 53.715 192.295 55.775 ;
        RECT 192.095 53.395 192.355 53.715 ;
        RECT 191.175 53.285 191.435 53.375 ;
        RECT 190.775 53.145 191.435 53.285 ;
        RECT 190.775 50.995 190.915 53.145 ;
        RECT 191.175 53.055 191.435 53.145 ;
        RECT 193.075 51.335 193.215 64.275 ;
        RECT 193.535 53.375 193.675 72.435 ;
        RECT 194.395 69.375 194.655 69.695 ;
        RECT 193.935 68.870 194.195 69.015 ;
        RECT 193.925 68.500 194.205 68.870 ;
        RECT 193.935 66.315 194.195 66.635 ;
        RECT 193.995 63.915 194.135 66.315 ;
        RECT 194.455 65.470 194.595 69.375 ;
        RECT 194.385 65.100 194.665 65.470 ;
        RECT 194.915 64.935 195.055 85.695 ;
        RECT 195.375 80.575 195.515 88.415 ;
        RECT 195.835 81.255 195.975 88.755 ;
        RECT 196.225 86.180 196.505 86.550 ;
        RECT 196.295 86.015 196.435 86.180 ;
        RECT 196.235 85.695 196.495 86.015 ;
        RECT 196.695 85.870 196.955 86.015 ;
        RECT 196.685 85.500 196.965 85.870 ;
        RECT 195.775 80.935 196.035 81.255 ;
        RECT 195.315 80.255 195.575 80.575 ;
        RECT 195.375 78.535 195.515 80.255 ;
        RECT 195.835 78.875 195.975 80.935 ;
        RECT 197.675 79.895 197.815 102.015 ;
        RECT 199.055 100.635 199.195 105.075 ;
        RECT 200.895 103.355 201.035 109.225 ;
        RECT 202.215 105.075 202.475 105.395 ;
        RECT 200.835 103.035 201.095 103.355 ;
        RECT 199.455 102.015 199.715 102.335 ;
        RECT 198.995 100.315 199.255 100.635 ;
        RECT 198.995 96.575 199.255 96.895 ;
        RECT 199.055 93.835 199.195 96.575 ;
        RECT 198.995 93.515 199.255 93.835 ;
        RECT 198.075 90.455 198.335 90.775 ;
        RECT 197.615 79.575 197.875 79.895 ;
        RECT 195.775 78.555 196.035 78.875 ;
        RECT 195.315 78.215 195.575 78.535 ;
        RECT 196.685 78.020 196.965 78.390 ;
        RECT 196.695 77.875 196.955 78.020 ;
        RECT 197.155 77.875 197.415 78.195 ;
        RECT 195.775 69.035 196.035 69.355 ;
        RECT 194.855 64.615 195.115 64.935 ;
        RECT 194.395 63.935 194.655 64.255 ;
        RECT 193.935 63.595 194.195 63.915 ;
        RECT 194.455 62.215 194.595 63.935 ;
        RECT 195.835 63.915 195.975 69.035 ;
        RECT 196.225 68.500 196.505 68.870 ;
        RECT 195.775 63.595 196.035 63.915 ;
        RECT 195.835 63.430 195.975 63.595 ;
        RECT 195.765 63.060 196.045 63.430 ;
        RECT 194.395 61.895 194.655 62.215 ;
        RECT 193.925 58.980 194.205 59.350 ;
        RECT 193.935 58.835 194.195 58.980 ;
        RECT 193.935 55.775 194.195 56.095 ;
        RECT 193.475 53.055 193.735 53.375 ;
        RECT 193.995 53.035 194.135 55.775 ;
        RECT 194.455 54.055 194.595 61.895 ;
        RECT 196.295 61.275 196.435 68.500 ;
        RECT 196.685 67.820 196.965 68.190 ;
        RECT 196.755 67.315 196.895 67.820 ;
        RECT 196.695 66.995 196.955 67.315 ;
        RECT 197.215 66.830 197.355 77.875 ;
        RECT 197.615 66.995 197.875 67.315 ;
        RECT 197.145 66.460 197.425 66.830 ;
        RECT 196.685 65.100 196.965 65.470 ;
        RECT 196.695 64.955 196.955 65.100 ;
        RECT 197.215 62.555 197.355 66.460 ;
        RECT 197.675 64.255 197.815 66.995 ;
        RECT 197.615 63.935 197.875 64.255 ;
        RECT 197.675 62.555 197.815 63.935 ;
        RECT 197.155 62.235 197.415 62.555 ;
        RECT 197.615 62.235 197.875 62.555 ;
        RECT 198.135 61.875 198.275 90.455 ;
        RECT 198.535 85.015 198.795 85.335 ;
        RECT 198.595 61.875 198.735 85.015 ;
        RECT 198.995 77.875 199.255 78.195 ;
        RECT 199.055 67.315 199.195 77.875 ;
        RECT 199.515 76.155 199.655 102.015 ;
        RECT 199.905 100.460 200.185 100.830 ;
        RECT 199.915 100.315 200.175 100.460 ;
        RECT 199.975 88.055 200.115 100.315 ;
        RECT 200.375 99.295 200.635 99.615 ;
        RECT 200.435 97.235 200.575 99.295 ;
        RECT 200.375 96.915 200.635 97.235 ;
        RECT 200.375 95.895 200.635 96.215 ;
        RECT 200.435 91.455 200.575 95.895 ;
        RECT 200.375 91.135 200.635 91.455 ;
        RECT 201.755 88.755 202.015 89.075 ;
        RECT 201.815 88.395 201.955 88.755 ;
        RECT 201.755 88.075 202.015 88.395 ;
        RECT 199.915 87.735 200.175 88.055 ;
        RECT 201.815 86.015 201.955 88.075 ;
        RECT 201.755 85.695 202.015 86.015 ;
        RECT 201.295 85.015 201.555 85.335 ;
        RECT 199.915 82.975 200.175 83.295 ;
        RECT 199.455 75.835 199.715 76.155 ;
        RECT 199.975 67.315 200.115 82.975 ;
        RECT 200.375 78.555 200.635 78.875 ;
        RECT 200.435 77.855 200.575 78.555 ;
        RECT 200.375 77.535 200.635 77.855 ;
        RECT 200.375 75.835 200.635 76.155 ;
        RECT 200.435 73.435 200.575 75.835 ;
        RECT 200.375 73.115 200.635 73.435 ;
        RECT 200.835 72.270 201.095 72.415 ;
        RECT 200.825 71.900 201.105 72.270 ;
        RECT 200.375 69.375 200.635 69.695 ;
        RECT 198.995 66.995 199.255 67.315 ;
        RECT 199.915 66.995 200.175 67.315 ;
        RECT 199.055 66.635 199.195 66.995 ;
        RECT 198.995 66.315 199.255 66.635 ;
        RECT 199.055 64.165 199.195 66.315 ;
        RECT 199.975 65.275 200.115 66.995 ;
        RECT 200.435 66.150 200.575 69.375 ;
        RECT 200.895 69.355 201.035 71.900 ;
        RECT 200.835 69.035 201.095 69.355 ;
        RECT 200.835 66.830 201.095 66.975 ;
        RECT 200.825 66.460 201.105 66.830 ;
        RECT 201.355 66.295 201.495 85.015 ;
        RECT 202.275 78.195 202.415 105.075 ;
        RECT 202.675 102.015 202.935 102.335 ;
        RECT 202.735 91.310 202.875 102.015 ;
        RECT 203.195 97.915 203.335 109.225 ;
        RECT 204.055 106.775 204.315 107.095 ;
        RECT 204.115 104.715 204.255 106.775 ;
        RECT 205.495 106.075 205.635 109.225 ;
        RECT 205.435 105.755 205.695 106.075 ;
        RECT 205.895 105.075 206.155 105.395 ;
        RECT 204.055 104.395 204.315 104.715 ;
        RECT 205.435 104.055 205.695 104.375 ;
        RECT 205.495 103.355 205.635 104.055 ;
        RECT 205.435 103.035 205.695 103.355 ;
        RECT 203.595 101.675 203.855 101.995 ;
        RECT 203.135 97.595 203.395 97.915 ;
        RECT 203.135 93.855 203.395 94.175 ;
        RECT 202.665 90.940 202.945 91.310 ;
        RECT 203.195 89.075 203.335 93.855 ;
        RECT 203.655 90.775 203.795 101.675 ;
        RECT 204.975 98.615 205.235 98.935 ;
        RECT 204.055 97.595 204.315 97.915 ;
        RECT 204.115 94.515 204.255 97.595 ;
        RECT 205.035 97.235 205.175 98.615 ;
        RECT 204.975 96.915 205.235 97.235 ;
        RECT 205.035 96.215 205.175 96.915 ;
        RECT 204.975 95.895 205.235 96.215 ;
        RECT 204.055 94.195 204.315 94.515 ;
        RECT 203.595 90.455 203.855 90.775 ;
        RECT 203.655 89.075 203.795 90.455 ;
        RECT 203.135 88.755 203.395 89.075 ;
        RECT 203.595 88.755 203.855 89.075 ;
        RECT 202.215 77.875 202.475 78.195 ;
        RECT 201.755 76.855 202.015 77.175 ;
        RECT 200.365 65.780 200.645 66.150 ;
        RECT 201.295 65.975 201.555 66.295 ;
        RECT 199.915 64.955 200.175 65.275 ;
        RECT 199.915 64.165 200.175 64.255 ;
        RECT 199.055 64.025 200.175 64.165 ;
        RECT 199.915 63.935 200.175 64.025 ;
        RECT 200.435 63.915 200.575 65.780 ;
        RECT 201.355 64.595 201.495 65.975 ;
        RECT 201.295 64.275 201.555 64.595 ;
        RECT 200.375 63.595 200.635 63.915 ;
        RECT 198.995 63.255 199.255 63.575 ;
        RECT 199.055 61.875 199.195 63.255 ;
        RECT 198.075 61.555 198.335 61.875 ;
        RECT 198.535 61.555 198.795 61.875 ;
        RECT 198.995 61.555 199.255 61.875 ;
        RECT 199.915 61.555 200.175 61.875 ;
        RECT 200.375 61.555 200.635 61.875 ;
        RECT 196.295 61.135 196.895 61.275 ;
        RECT 196.235 60.535 196.495 60.855 ;
        RECT 195.305 58.980 195.585 59.350 ;
        RECT 195.315 58.835 195.575 58.980 ;
        RECT 195.775 58.495 196.035 58.815 ;
        RECT 195.835 55.415 195.975 58.495 ;
        RECT 196.295 56.775 196.435 60.535 ;
        RECT 196.755 59.495 196.895 61.135 ;
        RECT 196.695 59.175 196.955 59.495 ;
        RECT 199.975 58.815 200.115 61.555 ;
        RECT 200.435 61.195 200.575 61.555 ;
        RECT 200.375 60.875 200.635 61.195 ;
        RECT 201.815 59.495 201.955 76.855 ;
        RECT 202.275 76.155 202.415 77.875 ;
        RECT 202.215 75.835 202.475 76.155 ;
        RECT 202.215 73.115 202.475 73.435 ;
        RECT 202.275 64.790 202.415 73.115 ;
        RECT 203.195 67.995 203.335 88.755 ;
        RECT 204.115 73.095 204.255 94.195 ;
        RECT 205.955 93.915 206.095 105.075 ;
        RECT 207.795 104.715 207.935 109.225 ;
        RECT 209.115 108.135 209.375 108.455 ;
        RECT 209.175 106.075 209.315 108.135 ;
        RECT 210.095 107.095 210.235 109.225 ;
        RECT 210.035 106.775 210.295 107.095 ;
        RECT 208.195 105.755 208.455 106.075 ;
        RECT 209.115 105.755 209.375 106.075 ;
        RECT 207.735 104.395 207.995 104.715 ;
        RECT 206.355 104.055 206.615 104.375 ;
        RECT 206.415 101.995 206.555 104.055 ;
        RECT 206.355 101.675 206.615 101.995 ;
        RECT 206.415 97.175 207.935 97.315 ;
        RECT 206.415 96.895 206.555 97.175 ;
        RECT 207.795 96.895 207.935 97.175 ;
        RECT 206.355 96.575 206.615 96.895 ;
        RECT 206.815 96.635 207.075 96.895 ;
        RECT 206.815 96.575 207.475 96.635 ;
        RECT 207.735 96.575 207.995 96.895 ;
        RECT 205.495 93.775 206.095 93.915 ;
        RECT 206.415 93.915 206.555 96.575 ;
        RECT 206.875 96.495 207.475 96.575 ;
        RECT 206.815 95.895 207.075 96.215 ;
        RECT 206.875 94.515 207.015 95.895 ;
        RECT 206.815 94.195 207.075 94.515 ;
        RECT 206.415 93.775 207.015 93.915 ;
        RECT 204.515 91.815 204.775 92.135 ;
        RECT 204.575 89.075 204.715 91.815 ;
        RECT 204.515 88.755 204.775 89.075 ;
        RECT 204.975 81.275 205.235 81.595 ;
        RECT 205.035 80.575 205.175 81.275 ;
        RECT 204.975 80.255 205.235 80.575 ;
        RECT 205.035 78.535 205.175 80.255 ;
        RECT 204.975 78.215 205.235 78.535 ;
        RECT 205.495 75.815 205.635 93.775 ;
        RECT 205.895 93.175 206.155 93.495 ;
        RECT 205.955 91.795 206.095 93.175 ;
        RECT 205.895 91.475 206.155 91.795 ;
        RECT 205.895 87.735 206.155 88.055 ;
        RECT 205.955 86.015 206.095 87.735 ;
        RECT 205.895 85.695 206.155 86.015 ;
        RECT 206.875 82.955 207.015 93.775 ;
        RECT 207.335 91.455 207.475 96.495 ;
        RECT 208.255 95.195 208.395 105.755 ;
        RECT 208.655 105.075 208.915 105.395 ;
        RECT 208.715 102.190 208.855 105.075 ;
        RECT 208.645 101.820 208.925 102.190 ;
        RECT 208.715 96.895 208.855 101.820 ;
        RECT 208.655 96.575 208.915 96.895 ;
        RECT 208.655 95.895 208.915 96.215 ;
        RECT 208.195 94.875 208.455 95.195 ;
        RECT 208.715 94.515 208.855 95.895 ;
        RECT 208.655 94.195 208.915 94.515 ;
        RECT 209.175 94.030 209.315 105.755 ;
        RECT 211.875 102.355 212.135 102.675 ;
        RECT 210.035 102.015 210.295 102.335 ;
        RECT 210.095 100.295 210.235 102.015 ;
        RECT 210.035 99.975 210.295 100.295 ;
        RECT 211.935 99.615 212.075 102.355 ;
        RECT 212.395 100.635 212.535 109.225 ;
        RECT 213.255 105.075 213.515 105.395 ;
        RECT 212.795 102.355 213.055 102.675 ;
        RECT 212.855 102.190 212.995 102.355 ;
        RECT 212.785 101.820 213.065 102.190 ;
        RECT 212.795 101.335 213.055 101.655 ;
        RECT 212.335 100.315 212.595 100.635 ;
        RECT 212.855 100.295 212.995 101.335 ;
        RECT 212.795 99.975 213.055 100.295 ;
        RECT 211.875 99.295 212.135 99.615 ;
        RECT 210.495 97.595 210.755 97.915 ;
        RECT 210.035 97.145 210.295 97.235 ;
        RECT 209.635 97.005 210.295 97.145 ;
        RECT 209.635 94.515 209.775 97.005 ;
        RECT 210.035 96.915 210.295 97.005 ;
        RECT 210.035 94.875 210.295 95.195 ;
        RECT 210.095 94.515 210.235 94.875 ;
        RECT 210.555 94.515 210.695 97.595 ;
        RECT 209.575 94.195 209.835 94.515 ;
        RECT 210.035 94.195 210.295 94.515 ;
        RECT 210.495 94.195 210.755 94.515 ;
        RECT 209.105 93.660 209.385 94.030 ;
        RECT 210.485 91.620 210.765 91.990 ;
        RECT 210.495 91.475 210.755 91.620 ;
        RECT 207.275 91.135 207.535 91.455 ;
        RECT 209.115 91.135 209.375 91.455 ;
        RECT 210.955 91.135 211.215 91.455 ;
        RECT 211.415 91.135 211.675 91.455 ;
        RECT 207.335 87.795 207.475 91.135 ;
        RECT 207.735 90.455 207.995 90.775 ;
        RECT 207.795 89.075 207.935 90.455 ;
        RECT 207.735 88.755 207.995 89.075 ;
        RECT 209.175 88.735 209.315 91.135 ;
        RECT 211.015 89.755 211.155 91.135 ;
        RECT 210.955 89.435 211.215 89.755 ;
        RECT 209.115 88.415 209.375 88.735 ;
        RECT 210.035 88.075 210.295 88.395 ;
        RECT 207.335 87.655 208.395 87.795 ;
        RECT 209.115 87.735 209.375 88.055 ;
        RECT 207.735 85.015 207.995 85.335 ;
        RECT 206.815 82.635 207.075 82.955 ;
        RECT 206.355 79.915 206.615 80.235 ;
        RECT 206.415 77.175 206.555 79.915 ;
        RECT 206.875 77.175 207.015 82.635 ;
        RECT 207.275 80.595 207.535 80.915 ;
        RECT 207.335 78.535 207.475 80.595 ;
        RECT 207.275 78.215 207.535 78.535 ;
        RECT 206.355 76.855 206.615 77.175 ;
        RECT 206.815 76.855 207.075 77.175 ;
        RECT 205.435 75.495 205.695 75.815 ;
        RECT 204.055 72.775 204.315 73.095 ;
        RECT 204.975 72.775 205.235 73.095 ;
        RECT 204.055 72.095 204.315 72.415 ;
        RECT 203.595 71.755 203.855 72.075 ;
        RECT 203.655 70.795 203.795 71.755 ;
        RECT 204.115 71.735 204.255 72.095 ;
        RECT 204.515 71.755 204.775 72.075 ;
        RECT 204.055 71.415 204.315 71.735 ;
        RECT 204.575 70.795 204.715 71.755 ;
        RECT 203.655 70.655 204.715 70.795 ;
        RECT 205.035 69.015 205.175 72.775 ;
        RECT 204.975 68.695 205.235 69.015 ;
        RECT 203.135 67.675 203.395 67.995 ;
        RECT 204.505 67.820 204.785 68.190 ;
        RECT 202.675 66.315 202.935 66.635 ;
        RECT 202.205 64.420 202.485 64.790 ;
        RECT 201.755 59.175 202.015 59.495 ;
        RECT 202.735 59.155 202.875 66.315 ;
        RECT 204.575 64.255 204.715 67.820 ;
        RECT 206.815 64.955 207.075 65.275 ;
        RECT 207.275 64.955 207.535 65.275 ;
        RECT 204.515 63.935 204.775 64.255 ;
        RECT 206.875 64.110 207.015 64.955 ;
        RECT 207.335 64.255 207.475 64.955 ;
        RECT 206.805 63.740 207.085 64.110 ;
        RECT 207.275 63.935 207.535 64.255 ;
        RECT 207.335 62.555 207.475 63.935 ;
        RECT 207.275 62.235 207.535 62.555 ;
        RECT 203.135 61.215 203.395 61.535 ;
        RECT 202.675 58.835 202.935 59.155 ;
        RECT 199.915 58.495 200.175 58.815 ;
        RECT 198.065 56.940 198.345 57.310 ;
        RECT 198.135 56.775 198.275 56.940 ;
        RECT 196.235 56.455 196.495 56.775 ;
        RECT 198.075 56.455 198.335 56.775 ;
        RECT 195.775 55.095 196.035 55.415 ;
        RECT 194.395 53.735 194.655 54.055 ;
        RECT 193.935 52.715 194.195 53.035 ;
        RECT 193.015 51.015 193.275 51.335 ;
        RECT 190.715 50.675 190.975 50.995 ;
        RECT 190.255 49.995 190.515 50.315 ;
        RECT 190.775 48.955 190.915 50.675 ;
        RECT 193.995 50.655 194.135 52.715 ;
        RECT 194.855 52.375 195.115 52.695 ;
        RECT 194.915 51.675 195.055 52.375 ;
        RECT 194.855 51.355 195.115 51.675 ;
        RECT 198.135 51.335 198.275 56.455 ;
        RECT 198.995 53.735 199.255 54.055 ;
        RECT 198.535 52.715 198.795 53.035 ;
        RECT 198.075 51.015 198.335 51.335 ;
        RECT 193.935 50.335 194.195 50.655 ;
        RECT 190.715 48.635 190.975 48.955 ;
        RECT 189.335 45.235 189.595 45.555 ;
        RECT 187.955 44.215 188.215 44.535 ;
        RECT 189.395 38.075 189.535 45.235 ;
        RECT 193.995 44.535 194.135 50.335 ;
        RECT 198.135 45.895 198.275 51.015 ;
        RECT 198.595 50.655 198.735 52.715 ;
        RECT 199.055 52.695 199.195 53.735 ;
        RECT 199.975 53.715 200.115 58.495 ;
        RECT 201.755 57.815 202.015 58.135 ;
        RECT 199.915 53.395 200.175 53.715 ;
        RECT 198.995 52.375 199.255 52.695 ;
        RECT 200.835 52.375 201.095 52.695 ;
        RECT 198.535 50.335 198.795 50.655 ;
        RECT 198.595 47.935 198.735 50.335 ;
        RECT 198.535 47.615 198.795 47.935 ;
        RECT 199.055 46.235 199.195 52.375 ;
        RECT 200.895 51.675 201.035 52.375 ;
        RECT 200.835 51.355 201.095 51.675 ;
        RECT 200.895 48.275 201.035 51.355 ;
        RECT 201.815 49.975 201.955 57.815 ;
        RECT 203.195 57.115 203.335 61.215 ;
        RECT 207.795 61.195 207.935 85.015 ;
        RECT 208.255 80.235 208.395 87.655 ;
        RECT 208.655 86.715 208.915 87.035 ;
        RECT 208.715 86.015 208.855 86.715 ;
        RECT 208.655 85.695 208.915 86.015 ;
        RECT 208.645 82.100 208.925 82.470 ;
        RECT 208.715 80.575 208.855 82.100 ;
        RECT 208.655 80.255 208.915 80.575 ;
        RECT 208.195 79.915 208.455 80.235 ;
        RECT 208.195 72.435 208.455 72.755 ;
        RECT 208.255 62.555 208.395 72.435 ;
        RECT 208.655 71.415 208.915 71.735 ;
        RECT 208.715 69.355 208.855 71.415 ;
        RECT 208.655 69.035 208.915 69.355 ;
        RECT 208.655 63.935 208.915 64.255 ;
        RECT 208.715 63.575 208.855 63.935 ;
        RECT 208.655 63.255 208.915 63.575 ;
        RECT 208.195 62.235 208.455 62.555 ;
        RECT 209.175 61.875 209.315 87.735 ;
        RECT 210.095 86.355 210.235 88.075 ;
        RECT 211.475 87.035 211.615 91.135 ;
        RECT 211.415 86.715 211.675 87.035 ;
        RECT 210.035 86.035 210.295 86.355 ;
        RECT 210.495 85.695 210.755 86.015 ;
        RECT 210.555 83.975 210.695 85.695 ;
        RECT 210.495 83.655 210.755 83.975 ;
        RECT 211.935 83.635 212.075 99.295 ;
        RECT 212.795 87.735 213.055 88.055 ;
        RECT 212.325 86.860 212.605 87.230 ;
        RECT 212.395 86.015 212.535 86.860 ;
        RECT 212.855 86.355 212.995 87.735 ;
        RECT 212.795 86.035 213.055 86.355 ;
        RECT 212.335 85.695 212.595 86.015 ;
        RECT 213.315 85.675 213.455 105.075 ;
        RECT 214.695 103.355 214.835 109.225 ;
        RECT 216.995 106.075 217.135 109.225 ;
        RECT 216.935 105.755 217.195 106.075 ;
        RECT 216.935 105.075 217.195 105.395 ;
        RECT 217.395 105.075 217.655 105.395 ;
        RECT 217.855 105.075 218.115 105.395 ;
        RECT 218.315 105.075 218.575 105.395 ;
        RECT 214.635 103.035 214.895 103.355 ;
        RECT 213.715 101.335 213.975 101.655 ;
        RECT 215.095 101.335 215.355 101.655 ;
        RECT 216.995 101.565 217.135 105.075 ;
        RECT 217.455 104.910 217.595 105.075 ;
        RECT 217.385 104.540 217.665 104.910 ;
        RECT 217.395 101.565 217.655 101.655 ;
        RECT 216.995 101.510 217.655 101.565 ;
        RECT 216.995 101.425 217.665 101.510 ;
        RECT 213.775 97.915 213.915 101.335 ;
        RECT 215.155 100.830 215.295 101.335 ;
        RECT 217.385 101.140 217.665 101.425 ;
        RECT 215.085 100.460 215.365 100.830 ;
        RECT 215.555 99.635 215.815 99.955 ;
        RECT 214.175 98.955 214.435 99.275 ;
        RECT 214.235 97.915 214.375 98.955 ;
        RECT 213.715 97.595 213.975 97.915 ;
        RECT 214.175 97.595 214.435 97.915 ;
        RECT 215.095 94.875 215.355 95.195 ;
        RECT 214.175 93.175 214.435 93.495 ;
        RECT 214.235 89.075 214.375 93.175 ;
        RECT 215.155 92.475 215.295 94.875 ;
        RECT 215.095 92.155 215.355 92.475 ;
        RECT 214.635 91.815 214.895 92.135 ;
        RECT 214.695 90.775 214.835 91.815 ;
        RECT 214.635 90.455 214.895 90.775 ;
        RECT 214.695 89.075 214.835 90.455 ;
        RECT 214.175 88.755 214.435 89.075 ;
        RECT 214.635 88.755 214.895 89.075 ;
        RECT 213.255 85.355 213.515 85.675 ;
        RECT 212.335 83.995 212.595 84.315 ;
        RECT 211.875 83.315 212.135 83.635 ;
        RECT 210.095 78.195 211.615 78.275 ;
        RECT 210.035 78.135 211.615 78.195 ;
        RECT 210.035 77.875 210.295 78.135 ;
        RECT 211.475 77.855 211.615 78.135 ;
        RECT 210.495 77.535 210.755 77.855 ;
        RECT 211.415 77.535 211.675 77.855 ;
        RECT 210.555 73.095 210.695 77.535 ;
        RECT 211.935 75.475 212.075 83.315 ;
        RECT 212.395 78.195 212.535 83.995 ;
        RECT 215.085 83.460 215.365 83.830 ;
        RECT 215.095 83.315 215.355 83.460 ;
        RECT 212.795 81.275 213.055 81.595 ;
        RECT 212.855 80.575 212.995 81.275 ;
        RECT 212.795 80.255 213.055 80.575 ;
        RECT 215.095 80.255 215.355 80.575 ;
        RECT 215.155 78.875 215.295 80.255 ;
        RECT 215.615 79.750 215.755 99.635 ;
        RECT 217.915 96.895 218.055 105.075 ;
        RECT 218.375 103.015 218.515 105.075 ;
        RECT 219.295 104.375 219.435 109.225 ;
        RECT 221.595 105.055 221.735 109.225 ;
        RECT 221.995 107.795 222.255 108.115 ;
        RECT 222.055 105.055 222.195 107.795 ;
        RECT 223.895 106.075 224.035 109.225 ;
        RECT 223.835 105.755 224.095 106.075 ;
        RECT 221.535 104.735 221.795 105.055 ;
        RECT 221.995 104.735 222.255 105.055 ;
        RECT 220.615 104.395 220.875 104.715 ;
        RECT 219.235 104.055 219.495 104.375 ;
        RECT 219.695 104.055 219.955 104.375 ;
        RECT 218.315 102.695 218.575 103.015 ;
        RECT 219.755 100.295 219.895 104.055 ;
        RECT 220.675 100.830 220.815 104.395 ;
        RECT 222.055 103.435 222.195 104.735 ;
        RECT 221.595 103.295 222.195 103.435 ;
        RECT 226.195 103.355 226.335 109.225 ;
        RECT 228.495 106.075 228.635 109.225 ;
        RECT 229.355 107.115 229.615 107.435 ;
        RECT 228.435 105.755 228.695 106.075 ;
        RECT 226.585 104.540 226.865 104.910 ;
        RECT 227.055 104.735 227.315 105.055 ;
        RECT 220.605 100.460 220.885 100.830 ;
        RECT 219.695 99.975 219.955 100.295 ;
        RECT 221.595 98.110 221.735 103.295 ;
        RECT 226.135 103.035 226.395 103.355 ;
        RECT 221.995 102.355 222.255 102.675 ;
        RECT 222.055 101.995 222.195 102.355 ;
        RECT 226.135 102.015 226.395 102.335 ;
        RECT 221.995 101.675 222.255 101.995 ;
        RECT 222.055 100.295 222.195 101.675 ;
        RECT 221.995 99.975 222.255 100.295 ;
        RECT 221.525 97.740 221.805 98.110 ;
        RECT 217.855 96.575 218.115 96.895 ;
        RECT 216.935 93.175 217.195 93.495 ;
        RECT 216.015 91.135 216.275 91.455 ;
        RECT 215.545 79.380 215.825 79.750 ;
        RECT 215.095 78.555 215.355 78.875 ;
        RECT 212.335 77.875 212.595 78.195 ;
        RECT 212.795 76.855 213.055 77.175 ;
        RECT 212.335 75.835 212.595 76.155 ;
        RECT 211.875 75.155 212.135 75.475 ;
        RECT 210.495 72.775 210.755 73.095 ;
        RECT 209.575 70.395 209.835 70.715 ;
        RECT 209.635 64.255 209.775 70.395 ;
        RECT 210.025 67.140 210.305 67.510 ;
        RECT 209.575 63.935 209.835 64.255 ;
        RECT 210.095 63.915 210.235 67.140 ;
        RECT 210.555 66.635 210.695 72.775 ;
        RECT 210.955 72.095 211.215 72.415 ;
        RECT 211.015 70.230 211.155 72.095 ;
        RECT 211.405 71.220 211.685 71.590 ;
        RECT 210.945 69.860 211.225 70.230 ;
        RECT 211.475 67.315 211.615 71.220 ;
        RECT 211.935 70.035 212.075 75.155 ;
        RECT 212.395 74.795 212.535 75.835 ;
        RECT 212.335 74.475 212.595 74.795 ;
        RECT 211.875 69.715 212.135 70.035 ;
        RECT 212.395 69.355 212.535 74.475 ;
        RECT 212.335 69.035 212.595 69.355 ;
        RECT 212.855 68.755 212.995 76.855 ;
        RECT 215.085 74.620 215.365 74.990 ;
        RECT 215.155 74.455 215.295 74.620 ;
        RECT 215.095 74.135 215.355 74.455 ;
        RECT 215.095 72.665 215.355 72.755 ;
        RECT 215.615 72.665 215.755 79.380 ;
        RECT 215.095 72.525 215.755 72.665 ;
        RECT 215.095 72.435 215.355 72.525 ;
        RECT 213.255 72.270 213.515 72.415 ;
        RECT 213.245 71.900 213.525 72.270 ;
        RECT 214.175 72.095 214.435 72.415 ;
        RECT 214.635 72.095 214.895 72.415 ;
        RECT 213.255 71.415 213.515 71.735 ;
        RECT 211.935 68.615 212.995 68.755 ;
        RECT 211.935 67.315 212.075 68.615 ;
        RECT 213.315 68.075 213.455 71.415 ;
        RECT 212.395 67.935 213.455 68.075 ;
        RECT 210.955 66.995 211.215 67.315 ;
        RECT 211.415 66.995 211.675 67.315 ;
        RECT 211.875 66.995 212.135 67.315 ;
        RECT 210.495 66.315 210.755 66.635 ;
        RECT 210.495 64.275 210.755 64.595 ;
        RECT 210.035 63.595 210.295 63.915 ;
        RECT 208.655 61.555 208.915 61.875 ;
        RECT 209.115 61.555 209.375 61.875 ;
        RECT 207.735 60.875 207.995 61.195 ;
        RECT 207.275 60.535 207.535 60.855 ;
        RECT 203.595 58.495 203.855 58.815 ;
        RECT 203.135 56.795 203.395 57.115 ;
        RECT 203.655 54.395 203.795 58.495 ;
        RECT 206.815 56.455 207.075 56.775 ;
        RECT 204.515 56.115 204.775 56.435 ;
        RECT 203.595 54.075 203.855 54.395 ;
        RECT 204.055 52.715 204.315 53.035 ;
        RECT 204.115 50.510 204.255 52.715 ;
        RECT 204.045 50.140 204.325 50.510 ;
        RECT 204.055 49.995 204.315 50.140 ;
        RECT 201.755 49.655 202.015 49.975 ;
        RECT 200.835 47.955 201.095 48.275 ;
        RECT 198.995 45.915 199.255 46.235 ;
        RECT 198.075 45.575 198.335 45.895 ;
        RECT 193.935 44.215 194.195 44.535 ;
        RECT 193.015 41.835 193.275 42.155 ;
        RECT 194.395 41.835 194.655 42.155 ;
        RECT 192.095 39.455 192.355 39.775 ;
        RECT 189.335 37.755 189.595 38.075 ;
        RECT 187.495 34.355 187.755 34.675 ;
        RECT 192.155 33.655 192.295 39.455 ;
        RECT 193.075 37.055 193.215 41.835 ;
        RECT 194.455 40.795 194.595 41.835 ;
        RECT 198.135 41.815 198.275 45.575 ;
        RECT 199.055 45.555 199.195 45.915 ;
        RECT 198.995 45.235 199.255 45.555 ;
        RECT 200.895 42.835 201.035 47.955 ;
        RECT 204.575 45.555 204.715 56.115 ;
        RECT 206.875 54.395 207.015 56.455 ;
        RECT 206.815 54.075 207.075 54.395 ;
        RECT 207.335 51.335 207.475 60.535 ;
        RECT 208.715 57.115 208.855 61.555 ;
        RECT 210.035 58.155 210.295 58.475 ;
        RECT 208.655 56.795 208.915 57.115 ;
        RECT 209.565 56.940 209.845 57.310 ;
        RECT 209.635 56.435 209.775 56.940 ;
        RECT 209.575 56.115 209.835 56.435 ;
        RECT 207.275 51.015 207.535 51.335 ;
        RECT 207.735 48.295 207.995 48.615 ;
        RECT 204.515 45.235 204.775 45.555 ;
        RECT 207.795 45.215 207.935 48.295 ;
        RECT 209.575 45.575 209.835 45.895 ;
        RECT 207.735 44.895 207.995 45.215 ;
        RECT 202.675 44.555 202.935 44.875 ;
        RECT 200.835 42.515 201.095 42.835 ;
        RECT 198.075 41.495 198.335 41.815 ;
        RECT 194.395 40.475 194.655 40.795 ;
        RECT 198.135 40.455 198.275 41.495 ;
        RECT 200.895 40.795 201.035 42.515 ;
        RECT 200.835 40.475 201.095 40.795 ;
        RECT 198.075 40.135 198.335 40.455 ;
        RECT 193.015 36.735 193.275 37.055 ;
        RECT 196.235 36.735 196.495 37.055 ;
        RECT 193.935 36.395 194.195 36.715 ;
        RECT 193.475 36.055 193.735 36.375 ;
        RECT 193.535 35.355 193.675 36.055 ;
        RECT 193.475 35.035 193.735 35.355 ;
        RECT 192.095 33.335 192.355 33.655 ;
        RECT 191.635 31.975 191.895 32.295 ;
        RECT 186.575 30.955 186.835 31.275 ;
        RECT 189.795 30.955 190.055 31.275 ;
        RECT 186.115 29.595 186.375 29.915 ;
        RECT 185.655 29.255 185.915 29.575 ;
        RECT 178.755 28.575 179.015 28.895 ;
        RECT 185.195 28.575 185.455 28.895 ;
        RECT 177.645 27.360 179.185 27.730 ;
        RECT 186.635 26.855 186.775 30.955 ;
        RECT 189.335 27.895 189.595 28.215 ;
        RECT 186.575 26.535 186.835 26.855 ;
        RECT 189.395 26.515 189.535 27.895 ;
        RECT 189.855 27.195 189.995 30.955 ;
        RECT 191.695 28.895 191.835 31.975 ;
        RECT 192.155 30.935 192.295 33.335 ;
        RECT 193.995 31.615 194.135 36.395 ;
        RECT 196.295 32.635 196.435 36.735 ;
        RECT 198.135 35.355 198.275 40.135 ;
        RECT 198.535 39.455 198.795 39.775 ;
        RECT 198.595 37.395 198.735 39.455 ;
        RECT 198.535 37.075 198.795 37.395 ;
        RECT 198.075 35.035 198.335 35.355 ;
        RECT 199.915 35.035 200.175 35.355 ;
        RECT 198.535 34.695 198.795 35.015 ;
        RECT 196.235 32.315 196.495 32.635 ;
        RECT 196.695 31.635 196.955 31.955 ;
        RECT 193.935 31.295 194.195 31.615 ;
        RECT 192.095 30.615 192.355 30.935 ;
        RECT 196.755 29.915 196.895 31.635 ;
        RECT 196.695 29.595 196.955 29.915 ;
        RECT 198.595 29.235 198.735 34.695 ;
        RECT 198.535 28.915 198.795 29.235 ;
        RECT 191.635 28.575 191.895 28.895 ;
        RECT 198.595 27.195 198.735 28.915 ;
        RECT 189.795 26.875 190.055 27.195 ;
        RECT 198.535 26.875 198.795 27.195 ;
        RECT 79.810 25.165 127.975 26.265 ;
        RECT 175.535 26.195 175.795 26.515 ;
        RECT 176.915 26.195 177.175 26.515 ;
        RECT 189.335 26.195 189.595 26.515 ;
        RECT 199.975 26.175 200.115 35.035 ;
        RECT 200.895 34.675 201.035 40.475 ;
        RECT 202.735 39.775 202.875 44.555 ;
        RECT 207.275 44.215 207.535 44.535 ;
        RECT 204.055 41.835 204.315 42.155 ;
        RECT 204.115 40.795 204.255 41.835 ;
        RECT 204.055 40.475 204.315 40.795 ;
        RECT 207.335 39.775 207.475 44.215 ;
        RECT 209.115 41.835 209.375 42.155 ;
        RECT 208.655 39.795 208.915 40.115 ;
        RECT 202.675 39.455 202.935 39.775 ;
        RECT 207.275 39.455 207.535 39.775 ;
        RECT 208.715 36.715 208.855 39.795 ;
        RECT 208.655 36.395 208.915 36.715 ;
        RECT 202.675 36.055 202.935 36.375 ;
        RECT 206.815 36.055 207.075 36.375 ;
        RECT 202.735 35.015 202.875 36.055 ;
        RECT 202.675 34.695 202.935 35.015 ;
        RECT 200.835 34.355 201.095 34.675 ;
        RECT 200.895 31.275 201.035 34.355 ;
        RECT 206.875 32.635 207.015 36.055 ;
        RECT 206.815 32.315 207.075 32.635 ;
        RECT 200.835 30.955 201.095 31.275 ;
        RECT 200.375 30.615 200.635 30.935 ;
        RECT 200.435 28.895 200.575 30.615 ;
        RECT 200.895 29.915 201.035 30.955 ;
        RECT 200.835 29.595 201.095 29.915 ;
        RECT 200.375 28.575 200.635 28.895 ;
        RECT 206.875 26.515 207.015 32.315 ;
        RECT 208.715 29.915 208.855 36.395 ;
        RECT 209.175 35.015 209.315 41.835 ;
        RECT 209.635 39.775 209.775 45.575 ;
        RECT 210.095 43.515 210.235 58.155 ;
        RECT 210.555 56.630 210.695 64.275 ;
        RECT 211.015 61.875 211.155 66.995 ;
        RECT 212.395 66.975 212.535 67.935 ;
        RECT 213.705 67.140 213.985 67.510 ;
        RECT 213.715 66.995 213.975 67.140 ;
        RECT 212.335 66.655 212.595 66.975 ;
        RECT 211.875 66.315 212.135 66.635 ;
        RECT 213.705 66.460 213.985 66.830 ;
        RECT 211.935 64.255 212.075 66.315 ;
        RECT 213.255 65.975 213.515 66.295 ;
        RECT 211.875 63.935 212.135 64.255 ;
        RECT 212.795 64.110 213.055 64.255 ;
        RECT 210.955 61.555 211.215 61.875 ;
        RECT 211.015 59.155 211.155 61.555 ;
        RECT 211.935 61.535 212.075 63.935 ;
        RECT 212.785 63.740 213.065 64.110 ;
        RECT 213.315 62.750 213.455 65.975 ;
        RECT 213.775 65.275 213.915 66.460 ;
        RECT 213.715 64.955 213.975 65.275 ;
        RECT 213.715 63.595 213.975 63.915 ;
        RECT 213.245 62.380 213.525 62.750 ;
        RECT 212.325 61.700 212.605 62.070 ;
        RECT 212.335 61.555 212.595 61.700 ;
        RECT 213.775 61.535 213.915 63.595 ;
        RECT 211.875 61.215 212.135 61.535 ;
        RECT 213.715 61.215 213.975 61.535 ;
        RECT 211.875 60.535 212.135 60.855 ;
        RECT 210.955 58.835 211.215 59.155 ;
        RECT 210.485 56.260 210.765 56.630 ;
        RECT 211.015 55.755 211.155 58.835 ;
        RECT 210.955 55.435 211.215 55.755 ;
        RECT 211.935 53.715 212.075 60.535 ;
        RECT 214.235 59.745 214.375 72.095 ;
        RECT 214.695 70.715 214.835 72.095 ;
        RECT 215.615 70.715 215.755 72.525 ;
        RECT 214.635 70.395 214.895 70.715 ;
        RECT 215.555 70.395 215.815 70.715 ;
        RECT 214.695 66.635 214.835 70.395 ;
        RECT 215.555 66.825 215.815 67.145 ;
        RECT 214.635 66.315 214.895 66.635 ;
        RECT 215.095 66.205 215.355 66.295 ;
        RECT 215.615 66.205 215.755 66.825 ;
        RECT 215.095 66.065 215.755 66.205 ;
        RECT 215.095 65.975 215.355 66.065 ;
        RECT 215.155 63.915 215.295 65.975 ;
        RECT 215.555 64.955 215.815 65.275 ;
        RECT 215.615 64.255 215.755 64.955 ;
        RECT 215.555 63.935 215.815 64.255 ;
        RECT 215.095 63.595 215.355 63.915 ;
        RECT 216.075 61.875 216.215 91.135 ;
        RECT 216.995 89.075 217.135 93.175 ;
        RECT 219.235 90.455 219.495 90.775 ;
        RECT 216.935 88.755 217.195 89.075 ;
        RECT 219.295 88.735 219.435 90.455 ;
        RECT 219.235 88.415 219.495 88.735 ;
        RECT 220.155 85.695 220.415 86.015 ;
        RECT 216.475 85.015 216.735 85.335 ;
        RECT 216.535 61.875 216.675 85.015 ;
        RECT 217.395 82.975 217.655 83.295 ;
        RECT 216.935 75.495 217.195 75.815 ;
        RECT 216.995 74.795 217.135 75.495 ;
        RECT 216.935 74.475 217.195 74.795 ;
        RECT 217.455 73.395 217.595 82.975 ;
        RECT 220.215 78.875 220.355 85.695 ;
        RECT 220.615 79.575 220.875 79.895 ;
        RECT 220.675 78.875 220.815 79.575 ;
        RECT 220.155 78.555 220.415 78.875 ;
        RECT 220.615 78.555 220.875 78.875 ;
        RECT 218.315 77.195 218.575 77.515 ;
        RECT 217.855 75.155 218.115 75.475 ;
        RECT 216.995 73.255 217.595 73.395 ;
        RECT 216.995 65.275 217.135 73.255 ;
        RECT 217.395 72.435 217.655 72.755 ;
        RECT 217.455 70.375 217.595 72.435 ;
        RECT 217.915 72.270 218.055 75.155 ;
        RECT 218.375 74.455 218.515 77.195 ;
        RECT 218.775 75.495 219.035 75.815 ;
        RECT 218.315 74.310 218.575 74.455 ;
        RECT 218.305 73.940 218.585 74.310 ;
        RECT 217.845 71.900 218.125 72.270 ;
        RECT 217.915 70.715 218.055 71.900 ;
        RECT 217.855 70.395 218.115 70.715 ;
        RECT 217.395 70.055 217.655 70.375 ;
        RECT 217.395 69.375 217.655 69.695 ;
        RECT 217.455 69.015 217.595 69.375 ;
        RECT 217.395 68.695 217.655 69.015 ;
        RECT 218.315 68.870 218.575 69.015 ;
        RECT 218.305 68.500 218.585 68.870 ;
        RECT 218.835 67.655 218.975 75.495 ;
        RECT 219.235 74.475 219.495 74.795 ;
        RECT 219.685 74.620 219.965 74.990 ;
        RECT 219.295 73.095 219.435 74.475 ;
        RECT 219.755 74.455 219.895 74.620 ;
        RECT 219.695 74.135 219.955 74.455 ;
        RECT 220.215 73.395 220.355 78.555 ;
        RECT 222.055 76.155 222.195 99.975 ;
        RECT 226.195 99.615 226.335 102.015 ;
        RECT 226.655 100.635 226.795 104.540 ;
        RECT 227.115 102.585 227.255 104.735 ;
        RECT 227.515 102.585 227.775 102.675 ;
        RECT 227.115 102.445 227.775 102.585 ;
        RECT 227.115 100.635 227.255 102.445 ;
        RECT 227.515 102.355 227.775 102.445 ;
        RECT 229.415 101.995 229.555 107.115 ;
        RECT 230.795 106.075 230.935 109.225 ;
        RECT 232.115 108.815 232.375 109.135 ;
        RECT 230.735 105.755 230.995 106.075 ;
        RECT 230.275 105.415 230.535 105.735 ;
        RECT 229.815 104.910 230.075 105.055 ;
        RECT 229.805 104.540 230.085 104.910 ;
        RECT 228.435 101.675 228.695 101.995 ;
        RECT 229.355 101.675 229.615 101.995 ;
        RECT 226.595 100.315 226.855 100.635 ;
        RECT 227.055 100.315 227.315 100.635 ;
        RECT 227.975 99.635 228.235 99.955 ;
        RECT 226.135 99.295 226.395 99.615 ;
        RECT 224.295 98.955 224.555 99.275 ;
        RECT 224.355 98.675 224.495 98.955 ;
        RECT 228.035 98.935 228.175 99.635 ;
        RECT 227.975 98.790 228.235 98.935 ;
        RECT 223.895 98.535 224.495 98.675 ;
        RECT 223.895 96.555 224.035 98.535 ;
        RECT 227.965 98.420 228.245 98.790 ;
        RECT 225.275 97.915 226.795 97.995 ;
        RECT 225.215 97.855 226.795 97.915 ;
        RECT 225.215 97.595 225.475 97.855 ;
        RECT 226.655 97.575 226.795 97.855 ;
        RECT 226.595 97.255 226.855 97.575 ;
        RECT 227.965 97.060 228.245 97.430 ;
        RECT 228.035 96.895 228.175 97.060 ;
        RECT 225.215 96.805 225.475 96.895 ;
        RECT 225.215 96.665 225.875 96.805 ;
        RECT 225.215 96.575 225.475 96.665 ;
        RECT 223.835 96.235 224.095 96.555 ;
        RECT 223.375 94.535 223.635 94.855 ;
        RECT 223.435 91.455 223.575 94.535 ;
        RECT 223.375 91.135 223.635 91.455 ;
        RECT 223.435 86.355 223.575 91.135 ;
        RECT 223.895 87.035 224.035 96.235 ;
        RECT 225.205 94.340 225.485 94.710 ;
        RECT 224.755 93.515 225.015 93.835 ;
        RECT 224.815 91.455 224.955 93.515 ;
        RECT 224.755 91.135 225.015 91.455 ;
        RECT 225.275 91.115 225.415 94.340 ;
        RECT 225.735 93.495 225.875 96.665 ;
        RECT 227.975 96.575 228.235 96.895 ;
        RECT 228.495 96.750 228.635 101.675 ;
        RECT 229.815 101.510 230.075 101.655 ;
        RECT 229.805 101.140 230.085 101.510 ;
        RECT 228.895 99.975 229.155 100.295 ;
        RECT 227.515 95.895 227.775 96.215 ;
        RECT 226.595 94.425 226.855 94.515 ;
        RECT 226.195 94.285 226.855 94.425 ;
        RECT 225.675 93.175 225.935 93.495 ;
        RECT 225.215 90.795 225.475 91.115 ;
        RECT 224.295 90.455 224.555 90.775 ;
        RECT 224.355 89.415 224.495 90.455 ;
        RECT 224.295 89.095 224.555 89.415 ;
        RECT 225.675 88.755 225.935 89.075 ;
        RECT 224.755 88.590 225.015 88.735 ;
        RECT 224.745 88.220 225.025 88.590 ;
        RECT 225.735 88.055 225.875 88.755 ;
        RECT 225.675 87.735 225.935 88.055 ;
        RECT 223.835 86.715 224.095 87.035 ;
        RECT 225.675 86.715 225.935 87.035 ;
        RECT 223.375 86.035 223.635 86.355 ;
        RECT 223.435 81.595 223.575 86.035 ;
        RECT 225.215 85.355 225.475 85.675 ;
        RECT 224.745 82.100 225.025 82.470 ;
        RECT 223.375 81.275 223.635 81.595 ;
        RECT 223.835 80.595 224.095 80.915 ;
        RECT 223.895 80.235 224.035 80.595 ;
        RECT 223.835 79.915 224.095 80.235 ;
        RECT 224.815 79.895 224.955 82.100 ;
        RECT 224.755 79.575 225.015 79.895 ;
        RECT 221.995 75.835 222.255 76.155 ;
        RECT 219.755 73.255 220.355 73.395 ;
        RECT 219.235 72.775 219.495 73.095 ;
        RECT 219.235 72.095 219.495 72.415 ;
        RECT 219.295 70.715 219.435 72.095 ;
        RECT 219.235 70.395 219.495 70.715 ;
        RECT 218.775 67.335 219.035 67.655 ;
        RECT 218.315 67.225 218.575 67.315 ;
        RECT 217.455 67.085 218.575 67.225 ;
        RECT 217.455 66.830 217.595 67.085 ;
        RECT 218.315 66.995 218.575 67.085 ;
        RECT 217.385 66.460 217.665 66.830 ;
        RECT 219.755 66.715 219.895 73.255 ;
        RECT 222.055 73.095 222.195 75.835 ;
        RECT 221.995 72.775 222.255 73.095 ;
        RECT 220.615 68.695 220.875 69.015 ;
        RECT 220.155 67.675 220.415 67.995 ;
        RECT 220.215 67.315 220.355 67.675 ;
        RECT 220.155 66.995 220.415 67.315 ;
        RECT 220.675 66.830 220.815 68.695 ;
        RECT 221.995 67.675 222.255 67.995 ;
        RECT 217.915 66.575 219.895 66.715 ;
        RECT 216.935 64.955 217.195 65.275 ;
        RECT 216.935 64.110 217.195 64.255 ;
        RECT 216.925 63.740 217.205 64.110 ;
        RECT 215.555 61.555 215.815 61.875 ;
        RECT 216.015 61.555 216.275 61.875 ;
        RECT 216.475 61.555 216.735 61.875 ;
        RECT 214.235 59.605 214.835 59.745 ;
        RECT 214.175 58.835 214.435 59.155 ;
        RECT 213.705 56.940 213.985 57.310 ;
        RECT 213.255 56.115 213.515 56.435 ;
        RECT 213.315 54.395 213.455 56.115 ;
        RECT 213.255 54.075 213.515 54.395 ;
        RECT 211.875 53.395 212.135 53.715 ;
        RECT 211.415 52.375 211.675 52.695 ;
        RECT 211.475 50.995 211.615 52.375 ;
        RECT 211.415 50.675 211.675 50.995 ;
        RECT 213.775 50.655 213.915 56.940 ;
        RECT 214.235 51.675 214.375 58.835 ;
        RECT 214.695 55.835 214.835 59.605 ;
        RECT 215.615 57.115 215.755 61.555 ;
        RECT 215.555 56.795 215.815 57.115 ;
        RECT 216.005 56.260 216.285 56.630 ;
        RECT 216.015 56.115 216.275 56.260 ;
        RECT 214.695 55.755 216.215 55.835 ;
        RECT 214.695 55.695 216.275 55.755 ;
        RECT 216.015 55.435 216.275 55.695 ;
        RECT 215.095 55.095 215.355 55.415 ;
        RECT 214.175 51.355 214.435 51.675 ;
        RECT 214.235 50.655 214.375 51.355 ;
        RECT 215.155 51.335 215.295 55.095 ;
        RECT 215.095 51.015 215.355 51.335 ;
        RECT 213.715 50.335 213.975 50.655 ;
        RECT 214.175 50.335 214.435 50.655 ;
        RECT 214.235 47.935 214.375 50.335 ;
        RECT 215.555 49.655 215.815 49.975 ;
        RECT 215.615 47.935 215.755 49.655 ;
        RECT 214.175 47.615 214.435 47.935 ;
        RECT 215.555 47.615 215.815 47.935 ;
        RECT 217.395 46.935 217.655 47.255 ;
        RECT 212.795 44.895 213.055 45.215 ;
        RECT 210.035 43.195 210.295 43.515 ;
        RECT 210.495 41.495 210.755 41.815 ;
        RECT 210.555 40.795 210.695 41.495 ;
        RECT 210.495 40.475 210.755 40.795 ;
        RECT 209.575 39.455 209.835 39.775 ;
        RECT 212.335 36.055 212.595 36.375 ;
        RECT 209.115 34.695 209.375 35.015 ;
        RECT 209.175 31.615 209.315 34.695 ;
        RECT 210.035 33.335 210.295 33.655 ;
        RECT 209.115 31.295 209.375 31.615 ;
        RECT 208.655 29.595 208.915 29.915 ;
        RECT 210.095 29.235 210.235 33.335 ;
        RECT 212.395 31.955 212.535 36.055 ;
        RECT 212.855 34.675 212.995 44.895 ;
        RECT 216.475 44.215 216.735 44.535 ;
        RECT 214.175 42.515 214.435 42.835 ;
        RECT 214.235 40.115 214.375 42.515 ;
        RECT 216.535 42.155 216.675 44.215 ;
        RECT 216.475 41.835 216.735 42.155 ;
        RECT 217.455 40.795 217.595 46.935 ;
        RECT 217.915 46.235 218.055 66.575 ;
        RECT 220.155 66.315 220.415 66.635 ;
        RECT 220.605 66.460 220.885 66.830 ;
        RECT 218.305 65.780 218.585 66.150 ;
        RECT 219.235 65.975 219.495 66.295 ;
        RECT 218.375 64.790 218.515 65.780 ;
        RECT 218.305 64.420 218.585 64.790 ;
        RECT 218.775 64.275 219.035 64.595 ;
        RECT 218.315 63.255 218.575 63.575 ;
        RECT 218.375 58.135 218.515 63.255 ;
        RECT 218.835 62.750 218.975 64.275 ;
        RECT 219.295 64.255 219.435 65.975 ;
        RECT 219.695 64.955 219.955 65.275 ;
        RECT 219.755 64.255 219.895 64.955 ;
        RECT 219.235 63.935 219.495 64.255 ;
        RECT 219.695 63.935 219.955 64.255 ;
        RECT 218.765 62.380 219.045 62.750 ;
        RECT 220.215 59.235 220.355 66.315 ;
        RECT 221.525 65.100 221.805 65.470 ;
        RECT 221.075 64.275 221.335 64.595 ;
        RECT 220.615 63.935 220.875 64.255 ;
        RECT 220.675 62.215 220.815 63.935 ;
        RECT 221.135 62.555 221.275 64.275 ;
        RECT 221.595 62.750 221.735 65.100 ;
        RECT 221.075 62.235 221.335 62.555 ;
        RECT 221.525 62.380 221.805 62.750 ;
        RECT 220.615 61.895 220.875 62.215 ;
        RECT 222.055 62.070 222.195 67.675 ;
        RECT 221.985 61.700 222.265 62.070 ;
        RECT 221.535 61.215 221.795 61.535 ;
        RECT 221.075 60.875 221.335 61.195 ;
        RECT 220.215 59.155 220.815 59.235 ;
        RECT 220.215 59.095 220.875 59.155 ;
        RECT 220.615 58.835 220.875 59.095 ;
        RECT 218.315 57.815 218.575 58.135 ;
        RECT 218.775 56.795 219.035 57.115 ;
        RECT 218.315 56.115 218.575 56.435 ;
        RECT 217.855 45.915 218.115 46.235 ;
        RECT 217.915 41.815 218.055 45.915 ;
        RECT 217.855 41.495 218.115 41.815 ;
        RECT 217.395 40.475 217.655 40.795 ;
        RECT 214.175 39.795 214.435 40.115 ;
        RECT 218.375 39.775 218.515 56.115 ;
        RECT 218.835 53.375 218.975 56.795 ;
        RECT 219.235 56.455 219.495 56.775 ;
        RECT 219.295 53.375 219.435 56.455 ;
        RECT 221.135 54.395 221.275 60.875 ;
        RECT 221.595 59.835 221.735 61.215 ;
        RECT 221.535 59.515 221.795 59.835 ;
        RECT 224.815 59.595 224.955 79.575 ;
        RECT 225.275 72.415 225.415 85.355 ;
        RECT 225.735 74.310 225.875 86.715 ;
        RECT 226.195 80.915 226.335 94.285 ;
        RECT 226.595 94.195 226.855 94.285 ;
        RECT 227.575 94.175 227.715 95.895 ;
        RECT 228.035 95.195 228.175 96.575 ;
        RECT 228.425 96.380 228.705 96.750 ;
        RECT 228.435 95.895 228.695 96.215 ;
        RECT 227.975 94.875 228.235 95.195 ;
        RECT 227.965 94.340 228.245 94.710 ;
        RECT 227.975 94.195 228.235 94.340 ;
        RECT 227.515 93.855 227.775 94.175 ;
        RECT 227.515 93.175 227.775 93.495 ;
        RECT 227.975 93.175 228.235 93.495 ;
        RECT 227.055 92.155 227.315 92.475 ;
        RECT 226.595 91.135 226.855 91.455 ;
        RECT 226.655 89.415 226.795 91.135 ;
        RECT 227.115 89.755 227.255 92.155 ;
        RECT 227.055 89.435 227.315 89.755 ;
        RECT 226.595 89.095 226.855 89.415 ;
        RECT 227.575 88.985 227.715 93.175 ;
        RECT 228.035 91.455 228.175 93.175 ;
        RECT 227.975 91.135 228.235 91.455 ;
        RECT 227.975 88.985 228.235 89.075 ;
        RECT 227.115 88.845 228.235 88.985 ;
        RECT 226.595 88.415 226.855 88.735 ;
        RECT 226.655 87.035 226.795 88.415 ;
        RECT 226.595 86.715 226.855 87.035 ;
        RECT 226.595 86.035 226.855 86.355 ;
        RECT 226.655 82.955 226.795 86.035 ;
        RECT 226.595 82.635 226.855 82.955 ;
        RECT 226.135 80.595 226.395 80.915 ;
        RECT 226.585 80.740 226.865 81.110 ;
        RECT 226.655 79.895 226.795 80.740 ;
        RECT 226.595 79.575 226.855 79.895 ;
        RECT 226.595 77.195 226.855 77.515 ;
        RECT 225.665 73.940 225.945 74.310 ;
        RECT 225.215 72.095 225.475 72.415 ;
        RECT 225.275 69.695 225.415 72.095 ;
        RECT 225.215 69.375 225.475 69.695 ;
        RECT 225.215 63.935 225.475 64.255 ;
        RECT 225.275 63.315 225.415 63.935 ;
        RECT 226.135 63.595 226.395 63.915 ;
        RECT 225.275 63.175 225.875 63.315 ;
        RECT 225.215 60.535 225.475 60.855 ;
        RECT 224.355 59.455 224.955 59.595 ;
        RECT 221.525 58.980 221.805 59.350 ;
        RECT 221.075 54.075 221.335 54.395 ;
        RECT 221.595 53.375 221.735 58.980 ;
        RECT 222.915 58.155 223.175 58.475 ;
        RECT 222.455 57.815 222.715 58.135 ;
        RECT 218.775 53.055 219.035 53.375 ;
        RECT 219.235 53.055 219.495 53.375 ;
        RECT 221.535 53.285 221.795 53.375 ;
        RECT 221.535 53.145 222.195 53.285 ;
        RECT 221.535 53.055 221.795 53.145 ;
        RECT 222.055 51.675 222.195 53.145 ;
        RECT 221.995 51.355 222.255 51.675 ;
        RECT 222.515 47.255 222.655 57.815 ;
        RECT 222.975 56.775 223.115 58.155 ;
        RECT 222.915 56.455 223.175 56.775 ;
        RECT 222.975 52.695 223.115 56.455 ;
        RECT 223.835 55.095 224.095 55.415 ;
        RECT 222.915 52.375 223.175 52.695 ;
        RECT 222.975 50.995 223.115 52.375 ;
        RECT 222.915 50.675 223.175 50.995 ;
        RECT 222.915 49.655 223.175 49.975 ;
        RECT 222.455 46.935 222.715 47.255 ;
        RECT 222.975 46.235 223.115 49.655 ;
        RECT 223.895 48.955 224.035 55.095 ;
        RECT 223.835 48.635 224.095 48.955 ;
        RECT 223.835 47.955 224.095 48.275 ;
        RECT 222.915 45.915 223.175 46.235 ;
        RECT 218.775 44.895 219.035 45.215 ;
        RECT 218.315 39.455 218.575 39.775 ;
        RECT 214.175 39.005 214.435 39.095 ;
        RECT 214.175 38.865 214.835 39.005 ;
        RECT 214.175 38.775 214.435 38.865 ;
        RECT 214.695 38.075 214.835 38.865 ;
        RECT 218.835 38.075 218.975 44.895 ;
        RECT 221.995 42.175 222.255 42.495 ;
        RECT 222.055 40.455 222.195 42.175 ;
        RECT 222.975 40.455 223.115 45.915 ;
        RECT 223.895 45.555 224.035 47.955 ;
        RECT 223.835 45.235 224.095 45.555 ;
        RECT 223.375 44.555 223.635 44.875 ;
        RECT 223.835 44.555 224.095 44.875 ;
        RECT 223.435 43.175 223.575 44.555 ;
        RECT 223.375 42.855 223.635 43.175 ;
        RECT 223.895 42.835 224.035 44.555 ;
        RECT 224.355 43.515 224.495 59.455 ;
        RECT 224.755 58.155 225.015 58.475 ;
        RECT 224.815 45.555 224.955 58.155 ;
        RECT 225.275 56.775 225.415 60.535 ;
        RECT 225.735 59.155 225.875 63.175 ;
        RECT 226.195 61.195 226.335 63.595 ;
        RECT 226.655 61.875 226.795 77.195 ;
        RECT 227.115 70.375 227.255 88.845 ;
        RECT 227.975 88.755 228.235 88.845 ;
        RECT 227.975 86.715 228.235 87.035 ;
        RECT 227.515 83.655 227.775 83.975 ;
        RECT 227.575 80.235 227.715 83.655 ;
        RECT 228.035 83.635 228.175 86.715 ;
        RECT 228.495 85.870 228.635 95.895 ;
        RECT 228.955 92.475 229.095 99.975 ;
        RECT 229.355 99.470 229.615 99.615 ;
        RECT 229.345 99.100 229.625 99.470 ;
        RECT 229.415 95.390 229.555 99.100 ;
        RECT 229.345 95.020 229.625 95.390 ;
        RECT 228.895 92.155 229.155 92.475 ;
        RECT 228.955 91.705 229.095 92.155 ;
        RECT 229.355 91.705 229.615 91.795 ;
        RECT 228.955 91.565 229.615 91.705 ;
        RECT 229.355 91.475 229.615 91.565 ;
        RECT 228.895 90.795 229.155 91.115 ;
        RECT 228.955 87.035 229.095 90.795 ;
        RECT 229.875 89.755 230.015 101.140 ;
        RECT 229.815 89.435 230.075 89.755 ;
        RECT 228.895 86.715 229.155 87.035 ;
        RECT 228.425 85.500 228.705 85.870 ;
        RECT 228.895 85.695 229.155 86.015 ;
        RECT 228.435 85.015 228.695 85.335 ;
        RECT 228.495 83.635 228.635 85.015 ;
        RECT 227.975 83.315 228.235 83.635 ;
        RECT 228.435 83.315 228.695 83.635 ;
        RECT 228.955 83.545 229.095 85.695 ;
        RECT 230.335 84.315 230.475 105.415 ;
        RECT 232.175 105.395 232.315 108.815 ;
        RECT 233.095 106.075 233.235 109.225 ;
        RECT 234.875 109.155 235.135 109.475 ;
        RECT 235.325 109.225 235.605 125.445 ;
        RECT 237.625 109.225 237.905 126.025 ;
        RECT 239.925 109.225 240.205 126.605 ;
        RECT 242.225 109.225 242.505 127.185 ;
        RECT 244.525 109.225 244.805 127.765 ;
        RECT 246.825 109.225 247.105 128.345 ;
        RECT 249.125 109.225 249.405 128.925 ;
        RECT 251.425 109.225 251.705 129.505 ;
        RECT 253.725 109.225 254.005 130.085 ;
        RECT 256.025 109.225 256.305 130.665 ;
        RECT 258.325 109.225 258.605 131.245 ;
        RECT 260.625 109.225 260.905 131.825 ;
        RECT 262.925 109.225 263.205 132.405 ;
        RECT 233.035 105.755 233.295 106.075 ;
        RECT 234.935 105.395 235.075 109.155 ;
        RECT 235.395 106.075 235.535 109.225 ;
        RECT 237.695 106.075 237.835 109.225 ;
        RECT 239.015 108.475 239.275 108.795 ;
        RECT 235.335 105.755 235.595 106.075 ;
        RECT 237.635 105.755 237.895 106.075 ;
        RECT 239.075 105.395 239.215 108.475 ;
        RECT 232.115 105.075 232.375 105.395 ;
        RECT 234.875 105.075 235.135 105.395 ;
        RECT 239.015 105.075 239.275 105.395 ;
        RECT 239.475 104.735 239.735 105.055 ;
        RECT 232.575 102.190 232.835 102.335 ;
        RECT 232.565 101.820 232.845 102.190 ;
        RECT 231.655 96.575 231.915 96.895 ;
        RECT 231.715 95.195 231.855 96.575 ;
        RECT 232.115 96.235 232.375 96.555 ;
        RECT 233.955 96.235 234.215 96.555 ;
        RECT 231.655 94.875 231.915 95.195 ;
        RECT 230.735 91.815 230.995 92.135 ;
        RECT 230.795 91.455 230.935 91.815 ;
        RECT 231.715 91.455 231.855 94.875 ;
        RECT 230.735 91.135 230.995 91.455 ;
        RECT 231.655 91.135 231.915 91.455 ;
        RECT 230.735 90.455 230.995 90.775 ;
        RECT 231.195 90.455 231.455 90.775 ;
        RECT 230.795 88.055 230.935 90.455 ;
        RECT 231.255 89.075 231.395 90.455 ;
        RECT 231.195 88.755 231.455 89.075 ;
        RECT 230.735 87.735 230.995 88.055 ;
        RECT 230.275 83.995 230.535 84.315 ;
        RECT 229.355 83.545 229.615 83.635 ;
        RECT 228.955 83.405 229.615 83.545 ;
        RECT 228.035 82.615 228.175 83.315 ;
        RECT 227.975 82.295 228.235 82.615 ;
        RECT 227.515 79.915 227.775 80.235 ;
        RECT 227.575 78.195 227.715 79.915 ;
        RECT 228.435 79.575 228.695 79.895 ;
        RECT 227.975 78.555 228.235 78.875 ;
        RECT 227.515 77.875 227.775 78.195 ;
        RECT 228.035 75.475 228.175 78.555 ;
        RECT 228.495 78.535 228.635 79.575 ;
        RECT 228.955 78.875 229.095 83.405 ;
        RECT 229.355 83.315 229.615 83.405 ;
        RECT 229.355 82.635 229.615 82.955 ;
        RECT 229.415 81.255 229.555 82.635 ;
        RECT 229.355 80.935 229.615 81.255 ;
        RECT 230.335 80.995 230.475 83.995 ;
        RECT 228.895 78.555 229.155 78.875 ;
        RECT 228.435 78.215 228.695 78.535 ;
        RECT 229.415 77.175 229.555 80.935 ;
        RECT 230.335 80.855 230.935 80.995 ;
        RECT 230.275 80.315 230.535 80.575 ;
        RECT 229.875 80.255 230.535 80.315 ;
        RECT 229.875 80.175 230.475 80.255 ;
        RECT 229.355 76.855 229.615 77.175 ;
        RECT 227.975 75.155 228.235 75.475 ;
        RECT 227.505 73.940 227.785 74.310 ;
        RECT 227.575 73.095 227.715 73.940 ;
        RECT 227.515 72.775 227.775 73.095 ;
        RECT 229.875 72.755 230.015 80.175 ;
        RECT 230.795 73.395 230.935 80.855 ;
        RECT 231.655 80.430 231.915 80.575 ;
        RECT 231.645 80.060 231.925 80.430 ;
        RECT 231.655 79.575 231.915 79.895 ;
        RECT 231.715 78.195 231.855 79.575 ;
        RECT 231.655 77.875 231.915 78.195 ;
        RECT 230.795 73.255 231.395 73.395 ;
        RECT 231.255 72.755 231.395 73.255 ;
        RECT 229.815 72.435 230.075 72.755 ;
        RECT 230.735 72.435 230.995 72.755 ;
        RECT 231.195 72.435 231.455 72.755 ;
        RECT 227.055 70.055 227.315 70.375 ;
        RECT 229.875 69.550 230.015 72.435 ;
        RECT 230.795 72.075 230.935 72.435 ;
        RECT 230.735 71.755 230.995 72.075 ;
        RECT 230.795 69.695 230.935 71.755 ;
        RECT 229.805 69.180 230.085 69.550 ;
        RECT 230.735 69.375 230.995 69.695 ;
        RECT 231.255 66.035 231.395 72.435 ;
        RECT 232.175 72.075 232.315 96.235 ;
        RECT 232.575 95.895 232.835 96.215 ;
        RECT 232.635 93.835 232.775 95.895 ;
        RECT 232.575 93.515 232.835 93.835 ;
        RECT 232.635 91.455 232.775 93.515 ;
        RECT 234.015 93.495 234.155 96.235 ;
        RECT 234.865 94.340 235.145 94.710 ;
        RECT 235.335 94.535 235.595 94.855 ;
        RECT 233.955 93.175 234.215 93.495 ;
        RECT 234.935 93.235 235.075 94.340 ;
        RECT 235.395 94.030 235.535 94.535 ;
        RECT 235.325 93.660 235.605 94.030 ;
        RECT 233.035 92.155 233.295 92.475 ;
        RECT 233.095 91.795 233.235 92.155 ;
        RECT 233.035 91.475 233.295 91.795 ;
        RECT 232.575 91.135 232.835 91.455 ;
        RECT 233.035 85.695 233.295 86.015 ;
        RECT 233.095 81.595 233.235 85.695 ;
        RECT 233.495 82.295 233.755 82.615 ;
        RECT 233.035 81.275 233.295 81.595 ;
        RECT 232.575 79.575 232.835 79.895 ;
        RECT 233.095 79.805 233.235 81.275 ;
        RECT 233.555 80.575 233.695 82.295 ;
        RECT 234.015 81.255 234.155 93.175 ;
        RECT 234.935 93.095 235.535 93.235 ;
        RECT 233.955 80.935 234.215 81.255 ;
        RECT 235.395 81.110 235.535 93.095 ;
        RECT 233.495 80.255 233.755 80.575 ;
        RECT 233.095 79.665 233.695 79.805 ;
        RECT 232.635 77.855 232.775 79.575 ;
        RECT 232.575 77.535 232.835 77.855 ;
        RECT 232.115 71.755 232.375 72.075 ;
        RECT 232.575 71.415 232.835 71.735 ;
        RECT 232.115 70.055 232.375 70.375 ;
        RECT 231.655 69.715 231.915 70.035 ;
        RECT 230.795 65.895 231.395 66.035 ;
        RECT 230.795 61.875 230.935 65.895 ;
        RECT 231.185 65.100 231.465 65.470 ;
        RECT 231.255 63.575 231.395 65.100 ;
        RECT 231.715 63.915 231.855 69.715 ;
        RECT 232.175 67.315 232.315 70.055 ;
        RECT 232.635 67.655 232.775 71.415 ;
        RECT 232.575 67.335 232.835 67.655 ;
        RECT 232.115 66.995 232.375 67.315 ;
        RECT 232.575 65.975 232.835 66.295 ;
        RECT 232.635 64.935 232.775 65.975 ;
        RECT 232.575 64.615 232.835 64.935 ;
        RECT 231.655 63.595 231.915 63.915 ;
        RECT 231.195 63.255 231.455 63.575 ;
        RECT 231.255 62.555 231.395 63.255 ;
        RECT 231.195 62.235 231.455 62.555 ;
        RECT 226.595 61.555 226.855 61.875 ;
        RECT 230.735 61.555 230.995 61.875 ;
        RECT 226.135 60.875 226.395 61.195 ;
        RECT 228.895 60.535 229.155 60.855 ;
        RECT 225.675 58.835 225.935 59.155 ;
        RECT 225.215 56.455 225.475 56.775 ;
        RECT 225.735 53.035 225.875 58.835 ;
        RECT 227.515 58.495 227.775 58.815 ;
        RECT 227.975 58.495 228.235 58.815 ;
        RECT 227.575 57.310 227.715 58.495 ;
        RECT 227.505 56.940 227.785 57.310 ;
        RECT 228.035 56.515 228.175 58.495 ;
        RECT 228.955 56.775 229.095 60.535 ;
        RECT 229.355 58.155 229.615 58.475 ;
        RECT 229.415 56.775 229.555 58.155 ;
        RECT 227.575 56.435 228.175 56.515 ;
        RECT 228.895 56.455 229.155 56.775 ;
        RECT 229.355 56.455 229.615 56.775 ;
        RECT 227.515 56.375 228.175 56.435 ;
        RECT 227.515 56.115 227.775 56.375 ;
        RECT 227.575 53.715 227.715 56.115 ;
        RECT 227.515 53.395 227.775 53.715 ;
        RECT 225.675 52.715 225.935 53.035 ;
        RECT 225.215 51.355 225.475 51.675 ;
        RECT 225.275 48.955 225.415 51.355 ;
        RECT 225.215 48.635 225.475 48.955 ;
        RECT 225.275 45.555 225.415 48.635 ;
        RECT 224.755 45.235 225.015 45.555 ;
        RECT 225.215 45.235 225.475 45.555 ;
        RECT 224.295 43.195 224.555 43.515 ;
        RECT 224.355 42.915 224.495 43.195 ;
        RECT 223.835 42.515 224.095 42.835 ;
        RECT 224.355 42.775 224.955 42.915 ;
        RECT 221.995 40.135 222.255 40.455 ;
        RECT 222.915 40.135 223.175 40.455 ;
        RECT 221.075 38.775 221.335 39.095 ;
        RECT 214.635 37.755 214.895 38.075 ;
        RECT 218.775 37.755 219.035 38.075 ;
        RECT 215.555 37.075 215.815 37.395 ;
        RECT 214.635 36.055 214.895 36.375 ;
        RECT 212.795 34.355 213.055 34.675 ;
        RECT 214.695 31.955 214.835 36.055 ;
        RECT 215.615 32.635 215.755 37.075 ;
        RECT 218.835 37.055 218.975 37.755 ;
        RECT 221.135 37.395 221.275 38.775 ;
        RECT 221.075 37.075 221.335 37.395 ;
        RECT 218.775 36.735 219.035 37.055 ;
        RECT 216.475 36.395 216.735 36.715 ;
        RECT 215.555 32.315 215.815 32.635 ;
        RECT 212.335 31.635 212.595 31.955 ;
        RECT 214.635 31.635 214.895 31.955 ;
        RECT 210.035 28.915 210.295 29.235 ;
        RECT 212.395 27.195 212.535 31.635 ;
        RECT 216.535 31.615 216.675 36.395 ;
        RECT 217.395 36.055 217.655 36.375 ;
        RECT 217.455 33.655 217.595 36.055 ;
        RECT 222.055 35.015 222.195 40.135 ;
        RECT 222.915 38.775 223.175 39.095 ;
        RECT 222.975 37.395 223.115 38.775 ;
        RECT 223.895 37.395 224.035 42.515 ;
        RECT 224.815 42.495 224.955 42.775 ;
        RECT 224.755 42.175 225.015 42.495 ;
        RECT 225.735 40.455 225.875 52.715 ;
        RECT 226.135 50.675 226.395 50.995 ;
        RECT 226.195 47.595 226.335 50.675 ;
        RECT 227.575 48.275 227.715 53.395 ;
        RECT 227.975 53.055 228.235 53.375 ;
        RECT 228.035 50.655 228.175 53.055 ;
        RECT 227.975 50.335 228.235 50.655 ;
        RECT 228.035 48.275 228.175 50.335 ;
        RECT 227.515 47.955 227.775 48.275 ;
        RECT 227.975 47.955 228.235 48.275 ;
        RECT 226.135 47.275 226.395 47.595 ;
        RECT 228.035 44.875 228.175 47.955 ;
        RECT 228.895 47.615 229.155 47.935 ;
        RECT 228.435 45.235 228.695 45.555 ;
        RECT 227.975 44.555 228.235 44.875 ;
        RECT 228.495 44.535 228.635 45.235 ;
        RECT 228.435 44.215 228.695 44.535 ;
        RECT 226.595 41.495 226.855 41.815 ;
        RECT 226.655 40.795 226.795 41.495 ;
        RECT 226.595 40.475 226.855 40.795 ;
        RECT 228.495 40.455 228.635 44.215 ;
        RECT 228.955 43.515 229.095 47.615 ;
        RECT 229.415 47.595 229.555 56.455 ;
        RECT 230.795 56.095 230.935 61.555 ;
        RECT 232.575 60.535 232.835 60.855 ;
        RECT 232.635 59.155 232.775 60.535 ;
        RECT 232.575 58.835 232.835 59.155 ;
        RECT 230.735 55.775 230.995 56.095 ;
        RECT 231.655 50.335 231.915 50.655 ;
        RECT 232.115 50.335 232.375 50.655 ;
        RECT 231.715 48.955 231.855 50.335 ;
        RECT 231.655 48.635 231.915 48.955 ;
        RECT 229.355 47.275 229.615 47.595 ;
        RECT 229.415 44.535 229.555 47.275 ;
        RECT 229.815 45.575 230.075 45.895 ;
        RECT 229.355 44.215 229.615 44.535 ;
        RECT 228.895 43.195 229.155 43.515 ;
        RECT 225.675 40.135 225.935 40.455 ;
        RECT 228.435 40.135 228.695 40.455 ;
        RECT 229.875 39.775 230.015 45.575 ;
        RECT 232.175 45.215 232.315 50.335 ;
        RECT 232.115 44.895 232.375 45.215 ;
        RECT 232.575 44.215 232.835 44.535 ;
        RECT 232.115 41.495 232.375 41.815 ;
        RECT 232.175 40.795 232.315 41.495 ;
        RECT 232.115 40.475 232.375 40.795 ;
        RECT 227.975 39.455 228.235 39.775 ;
        RECT 229.815 39.455 230.075 39.775 ;
        RECT 225.675 38.775 225.935 39.095 ;
        RECT 222.915 37.075 223.175 37.395 ;
        RECT 223.835 37.075 224.095 37.395 ;
        RECT 221.995 34.695 222.255 35.015 ;
        RECT 223.895 34.335 224.035 37.075 ;
        RECT 225.735 37.055 225.875 38.775 ;
        RECT 225.675 36.735 225.935 37.055 ;
        RECT 225.675 36.055 225.935 36.375 ;
        RECT 225.735 35.015 225.875 36.055 ;
        RECT 225.675 34.695 225.935 35.015 ;
        RECT 222.455 34.015 222.715 34.335 ;
        RECT 223.835 34.015 224.095 34.335 ;
        RECT 217.395 33.335 217.655 33.655 ;
        RECT 219.235 33.335 219.495 33.655 ;
        RECT 219.295 31.615 219.435 33.335 ;
        RECT 222.515 32.635 222.655 34.015 ;
        RECT 222.455 32.315 222.715 32.635 ;
        RECT 223.895 31.955 224.035 34.015 ;
        RECT 223.835 31.635 224.095 31.955 ;
        RECT 228.035 31.615 228.175 39.455 ;
        RECT 230.275 38.775 230.535 39.095 ;
        RECT 230.335 37.395 230.475 38.775 ;
        RECT 230.275 37.075 230.535 37.395 ;
        RECT 232.635 34.675 232.775 44.215 ;
        RECT 233.555 42.915 233.695 79.665 ;
        RECT 234.015 78.535 234.155 80.935 ;
        RECT 235.325 80.740 235.605 81.110 ;
        RECT 235.395 80.575 235.535 80.740 ;
        RECT 239.535 80.575 239.675 104.735 ;
        RECT 239.995 103.435 240.135 109.225 ;
        RECT 240.855 107.795 241.115 108.115 ;
        RECT 240.915 105.395 241.055 107.795 ;
        RECT 242.295 106.075 242.435 109.225 ;
        RECT 244.595 107.095 244.735 109.225 ;
        RECT 244.535 106.775 244.795 107.095 ;
        RECT 242.235 105.755 242.495 106.075 ;
        RECT 240.855 105.075 241.115 105.395 ;
        RECT 245.915 105.075 246.175 105.395 ;
        RECT 239.995 103.355 240.595 103.435 ;
        RECT 239.995 103.295 240.655 103.355 ;
        RECT 240.395 103.035 240.655 103.295 ;
        RECT 240.915 96.750 241.055 105.075 ;
        RECT 242.695 104.395 242.955 104.715 ;
        RECT 241.315 104.055 241.575 104.375 ;
        RECT 241.375 100.295 241.515 104.055 ;
        RECT 242.755 101.655 242.895 104.395 ;
        RECT 245.975 103.015 246.115 105.075 ;
        RECT 245.915 102.695 246.175 103.015 ;
        RECT 242.695 101.335 242.955 101.655 ;
        RECT 241.315 99.975 241.575 100.295 ;
        RECT 242.695 97.255 242.955 97.575 ;
        RECT 240.845 96.380 241.125 96.750 ;
        RECT 241.775 96.575 242.035 96.895 ;
        RECT 241.315 96.235 241.575 96.555 ;
        RECT 241.375 94.710 241.515 96.235 ;
        RECT 241.305 94.340 241.585 94.710 ;
        RECT 241.835 93.495 241.975 96.575 ;
        RECT 242.755 94.855 242.895 97.255 ;
        RECT 243.605 97.060 243.885 97.430 ;
        RECT 244.535 97.255 244.795 97.575 ;
        RECT 243.675 96.895 243.815 97.060 ;
        RECT 243.615 96.575 243.875 96.895 ;
        RECT 242.695 94.535 242.955 94.855 ;
        RECT 242.695 93.855 242.955 94.175 ;
        RECT 241.775 93.175 242.035 93.495 ;
        RECT 240.855 91.135 241.115 91.455 ;
        RECT 240.395 86.715 240.655 87.035 ;
        RECT 240.455 81.255 240.595 86.715 ;
        RECT 240.395 80.935 240.655 81.255 ;
        RECT 240.915 80.995 241.055 91.135 ;
        RECT 242.755 87.035 242.895 93.855 ;
        RECT 243.155 90.795 243.415 91.115 ;
        RECT 243.615 90.795 243.875 91.115 ;
        RECT 242.695 86.715 242.955 87.035 ;
        RECT 241.315 85.355 241.575 85.675 ;
        RECT 241.375 82.615 241.515 85.355 ;
        RECT 242.695 83.655 242.955 83.975 ;
        RECT 242.755 83.150 242.895 83.655 ;
        RECT 242.685 82.780 242.965 83.150 ;
        RECT 241.315 82.295 241.575 82.615 ;
        RECT 242.235 82.295 242.495 82.615 ;
        RECT 243.215 82.355 243.355 90.795 ;
        RECT 243.675 90.630 243.815 90.795 ;
        RECT 243.605 90.260 243.885 90.630 ;
        RECT 243.615 87.735 243.875 88.055 ;
        RECT 243.675 86.550 243.815 87.735 ;
        RECT 244.595 87.230 244.735 97.255 ;
        RECT 245.975 94.175 246.115 102.695 ;
        RECT 246.375 101.675 246.635 101.995 ;
        RECT 246.435 100.295 246.575 101.675 ;
        RECT 246.375 99.975 246.635 100.295 ;
        RECT 246.895 99.275 247.035 109.225 ;
        RECT 248.675 107.795 248.935 108.115 ;
        RECT 248.735 105.395 248.875 107.795 ;
        RECT 249.195 106.075 249.335 109.225 ;
        RECT 249.135 105.755 249.395 106.075 ;
        RECT 248.675 105.075 248.935 105.395 ;
        RECT 247.755 104.735 248.015 105.055 ;
        RECT 247.815 102.335 247.955 104.735 ;
        RECT 251.495 104.715 251.635 109.225 ;
        RECT 253.275 108.815 253.535 109.135 ;
        RECT 252.815 107.455 253.075 107.775 ;
        RECT 252.875 105.055 253.015 107.455 ;
        RECT 252.815 104.735 253.075 105.055 ;
        RECT 249.135 104.395 249.395 104.715 ;
        RECT 251.435 104.395 251.695 104.715 ;
        RECT 248.675 104.055 248.935 104.375 ;
        RECT 248.735 102.675 248.875 104.055 ;
        RECT 249.195 102.675 249.335 104.395 ;
        RECT 248.675 102.355 248.935 102.675 ;
        RECT 249.135 102.355 249.395 102.675 ;
        RECT 247.755 102.015 248.015 102.335 ;
        RECT 246.835 98.955 247.095 99.275 ;
        RECT 247.815 98.935 247.955 102.015 ;
        RECT 248.215 101.335 248.475 101.655 ;
        RECT 251.895 101.335 252.155 101.655 ;
        RECT 247.755 98.615 248.015 98.935 ;
        RECT 247.295 97.595 247.555 97.915 ;
        RECT 246.835 96.575 247.095 96.895 ;
        RECT 246.375 95.895 246.635 96.215 ;
        RECT 246.895 96.070 247.035 96.575 ;
        RECT 244.995 93.855 245.255 94.175 ;
        RECT 245.915 93.855 246.175 94.175 ;
        RECT 245.055 89.075 245.195 93.855 ;
        RECT 245.915 93.350 246.175 93.495 ;
        RECT 245.905 92.980 246.185 93.350 ;
        RECT 245.455 91.815 245.715 92.135 ;
        RECT 244.995 88.755 245.255 89.075 ;
        RECT 245.515 88.735 245.655 91.815 ;
        RECT 245.975 91.455 246.115 92.980 ;
        RECT 245.915 91.135 246.175 91.455 ;
        RECT 246.435 89.075 246.575 95.895 ;
        RECT 246.825 95.700 247.105 96.070 ;
        RECT 247.355 94.515 247.495 97.595 ;
        RECT 247.295 94.195 247.555 94.515 ;
        RECT 247.295 93.515 247.555 93.835 ;
        RECT 247.355 90.775 247.495 93.515 ;
        RECT 247.815 91.455 247.955 98.615 ;
        RECT 248.275 98.110 248.415 101.335 ;
        RECT 251.955 100.295 252.095 101.335 ;
        RECT 251.895 99.975 252.155 100.295 ;
        RECT 249.135 98.615 249.395 98.935 ;
        RECT 248.205 97.740 248.485 98.110 ;
        RECT 249.195 97.575 249.335 98.615 ;
        RECT 249.135 97.255 249.395 97.575 ;
        RECT 248.275 96.555 249.795 96.635 ;
        RECT 250.055 96.575 250.315 96.895 ;
        RECT 248.215 96.495 249.795 96.555 ;
        RECT 248.215 96.235 248.475 96.495 ;
        RECT 248.675 95.895 248.935 96.215 ;
        RECT 248.735 94.855 248.875 95.895 ;
        RECT 249.655 95.105 249.795 96.495 ;
        RECT 250.115 96.070 250.255 96.575 ;
        RECT 251.895 96.235 252.155 96.555 ;
        RECT 250.045 95.700 250.325 96.070 ;
        RECT 250.515 95.105 250.775 95.195 ;
        RECT 249.655 94.965 250.775 95.105 ;
        RECT 250.515 94.875 250.775 94.965 ;
        RECT 248.675 94.535 248.935 94.855 ;
        RECT 249.125 94.340 249.405 94.710 ;
        RECT 251.955 94.515 252.095 96.235 ;
        RECT 249.135 94.195 249.395 94.340 ;
        RECT 251.435 94.195 251.695 94.515 ;
        RECT 251.895 94.195 252.155 94.515 ;
        RECT 252.355 94.195 252.615 94.515 ;
        RECT 252.805 94.340 253.085 94.710 ;
        RECT 252.815 94.195 253.075 94.340 ;
        RECT 248.675 93.855 248.935 94.175 ;
        RECT 248.215 93.175 248.475 93.495 ;
        RECT 248.275 91.455 248.415 93.175 ;
        RECT 247.755 91.135 248.015 91.455 ;
        RECT 248.215 91.135 248.475 91.455 ;
        RECT 247.295 90.455 247.555 90.775 ;
        RECT 247.755 90.455 248.015 90.775 ;
        RECT 246.375 88.755 246.635 89.075 ;
        RECT 245.455 88.415 245.715 88.735 ;
        RECT 246.835 88.590 247.095 88.735 ;
        RECT 246.825 88.220 247.105 88.590 ;
        RECT 247.295 87.735 247.555 88.055 ;
        RECT 244.525 86.860 244.805 87.230 ;
        RECT 243.605 86.180 243.885 86.550 ;
        RECT 244.535 86.375 244.795 86.695 ;
        RECT 244.595 83.975 244.735 86.375 ;
        RECT 244.995 85.015 245.255 85.335 ;
        RECT 244.535 83.715 244.795 83.975 ;
        RECT 244.135 83.655 244.795 83.715 ;
        RECT 243.615 83.315 243.875 83.635 ;
        RECT 244.135 83.575 244.735 83.655 ;
        RECT 245.055 83.635 245.195 85.015 ;
        RECT 247.355 83.635 247.495 87.735 ;
        RECT 247.815 86.695 247.955 90.455 ;
        RECT 247.755 86.375 248.015 86.695 ;
        RECT 247.755 85.870 248.015 86.015 ;
        RECT 247.745 85.500 248.025 85.870 ;
        RECT 248.275 83.975 248.415 91.135 ;
        RECT 248.735 91.115 248.875 93.855 ;
        RECT 250.515 93.175 250.775 93.495 ;
        RECT 250.975 93.175 251.235 93.495 ;
        RECT 251.495 93.350 251.635 94.195 ;
        RECT 250.575 91.990 250.715 93.175 ;
        RECT 251.035 92.475 251.175 93.175 ;
        RECT 251.425 92.980 251.705 93.350 ;
        RECT 250.975 92.155 251.235 92.475 ;
        RECT 250.505 91.620 250.785 91.990 ;
        RECT 248.675 90.795 248.935 91.115 ;
        RECT 250.515 88.755 250.775 89.075 ;
        RECT 250.575 87.035 250.715 88.755 ;
        RECT 251.495 88.055 251.635 92.980 ;
        RECT 251.435 87.735 251.695 88.055 ;
        RECT 250.515 86.715 250.775 87.035 ;
        RECT 252.415 86.695 252.555 94.195 ;
        RECT 252.875 88.395 253.015 94.195 ;
        RECT 252.815 88.075 253.075 88.395 ;
        RECT 252.355 86.375 252.615 86.695 ;
        RECT 248.675 86.035 248.935 86.355 ;
        RECT 248.215 83.655 248.475 83.975 ;
        RECT 248.735 83.635 248.875 86.035 ;
        RECT 249.135 85.695 249.395 86.015 ;
        RECT 242.295 81.595 242.435 82.295 ;
        RECT 242.755 82.215 243.355 82.355 ;
        RECT 242.235 81.275 242.495 81.595 ;
        RECT 240.455 80.575 240.595 80.935 ;
        RECT 240.915 80.855 241.515 80.995 ;
        RECT 234.415 80.315 234.675 80.575 ;
        RECT 234.415 80.255 235.075 80.315 ;
        RECT 235.335 80.255 235.595 80.575 ;
        RECT 239.475 80.255 239.735 80.575 ;
        RECT 240.395 80.255 240.655 80.575 ;
        RECT 240.855 80.255 241.115 80.575 ;
        RECT 234.475 80.175 235.075 80.255 ;
        RECT 233.955 78.215 234.215 78.535 ;
        RECT 234.935 73.395 235.075 80.175 ;
        RECT 238.555 74.815 238.815 75.135 ;
        RECT 234.935 73.255 235.535 73.395 ;
        RECT 234.415 72.435 234.675 72.755 ;
        RECT 234.475 70.035 234.615 72.435 ;
        RECT 234.415 69.715 234.675 70.035 ;
        RECT 234.865 69.860 235.145 70.230 ;
        RECT 234.935 66.830 235.075 69.860 ;
        RECT 235.395 69.015 235.535 73.255 ;
        RECT 236.255 69.435 236.515 69.695 ;
        RECT 236.255 69.375 236.915 69.435 ;
        RECT 236.315 69.295 236.915 69.375 ;
        RECT 235.335 68.870 235.595 69.015 ;
        RECT 235.325 68.500 235.605 68.870 ;
        RECT 236.255 68.695 236.515 69.015 ;
        RECT 236.315 66.975 236.455 68.695 ;
        RECT 234.865 66.460 235.145 66.830 ;
        RECT 235.795 66.655 236.055 66.975 ;
        RECT 236.255 66.655 236.515 66.975 ;
        RECT 234.935 61.875 235.075 66.460 ;
        RECT 235.855 66.150 235.995 66.655 ;
        RECT 235.785 65.780 236.065 66.150 ;
        RECT 236.775 61.875 236.915 69.295 ;
        RECT 234.875 61.555 235.135 61.875 ;
        RECT 236.715 61.555 236.975 61.875 ;
        RECT 238.095 55.775 238.355 56.095 ;
        RECT 238.155 54.395 238.295 55.775 ;
        RECT 238.095 54.075 238.355 54.395 ;
        RECT 237.175 50.675 237.435 50.995 ;
        RECT 237.235 45.555 237.375 50.675 ;
        RECT 237.175 45.465 237.435 45.555 ;
        RECT 236.775 45.325 237.435 45.465 ;
        RECT 235.335 44.895 235.595 45.215 ;
        RECT 233.095 42.775 233.695 42.915 ;
        RECT 233.095 40.115 233.235 42.775 ;
        RECT 235.395 42.495 235.535 44.895 ;
        RECT 236.255 42.745 236.515 42.835 ;
        RECT 236.775 42.745 236.915 45.325 ;
        RECT 237.175 45.235 237.435 45.325 ;
        RECT 236.255 42.605 236.915 42.745 ;
        RECT 236.255 42.515 236.515 42.605 ;
        RECT 233.495 42.175 233.755 42.495 ;
        RECT 235.335 42.175 235.595 42.495 ;
        RECT 233.035 39.795 233.295 40.115 ;
        RECT 233.095 38.075 233.235 39.795 ;
        RECT 233.035 37.755 233.295 38.075 ;
        RECT 233.555 35.355 233.695 42.175 ;
        RECT 236.775 36.715 236.915 42.605 ;
        RECT 237.175 42.175 237.435 42.495 ;
        RECT 237.235 40.795 237.375 42.175 ;
        RECT 238.615 41.815 238.755 74.815 ;
        RECT 239.015 69.375 239.275 69.695 ;
        RECT 239.075 66.150 239.215 69.375 ;
        RECT 239.005 65.780 239.285 66.150 ;
        RECT 239.075 62.070 239.215 65.780 ;
        RECT 239.535 62.555 239.675 80.255 ;
        RECT 240.915 73.395 241.055 80.255 ;
        RECT 241.375 74.795 241.515 80.855 ;
        RECT 241.765 80.740 242.045 81.110 ;
        RECT 241.835 80.575 241.975 80.740 ;
        RECT 241.775 80.255 242.035 80.575 ;
        RECT 242.235 77.875 242.495 78.195 ;
        RECT 241.315 74.475 241.575 74.795 ;
        RECT 240.455 73.255 241.055 73.395 ;
        RECT 240.455 69.695 240.595 73.255 ;
        RECT 241.775 72.950 242.035 73.095 ;
        RECT 240.855 72.435 241.115 72.755 ;
        RECT 241.765 72.580 242.045 72.950 ;
        RECT 240.915 70.910 241.055 72.435 ;
        RECT 241.775 71.755 242.035 72.075 ;
        RECT 241.315 71.415 241.575 71.735 ;
        RECT 240.845 70.540 241.125 70.910 ;
        RECT 240.395 69.375 240.655 69.695 ;
        RECT 239.935 68.695 240.195 69.015 ;
        RECT 240.395 68.695 240.655 69.015 ;
        RECT 239.475 62.235 239.735 62.555 ;
        RECT 239.005 61.700 239.285 62.070 ;
        RECT 239.535 59.835 239.675 62.235 ;
        RECT 239.475 59.515 239.735 59.835 ;
        RECT 239.995 59.350 240.135 68.695 ;
        RECT 240.455 67.995 240.595 68.695 ;
        RECT 240.395 67.675 240.655 67.995 ;
        RECT 240.855 67.675 241.115 67.995 ;
        RECT 240.915 67.315 241.055 67.675 ;
        RECT 241.375 67.315 241.515 71.415 ;
        RECT 240.855 66.995 241.115 67.315 ;
        RECT 241.315 66.995 241.575 67.315 ;
        RECT 241.315 66.315 241.575 66.635 ;
        RECT 241.375 65.275 241.515 66.315 ;
        RECT 241.835 66.295 241.975 71.755 ;
        RECT 242.295 66.715 242.435 77.875 ;
        RECT 242.755 67.225 242.895 82.215 ;
        RECT 243.675 81.595 243.815 83.315 ;
        RECT 243.615 81.275 243.875 81.595 ;
        RECT 244.135 80.575 244.275 83.575 ;
        RECT 244.995 83.315 245.255 83.635 ;
        RECT 246.375 83.315 246.635 83.635 ;
        RECT 247.295 83.315 247.555 83.635 ;
        RECT 248.675 83.315 248.935 83.635 ;
        RECT 246.435 80.915 246.575 83.315 ;
        RECT 247.355 83.035 247.495 83.315 ;
        RECT 246.895 82.895 247.495 83.035 ;
        RECT 247.755 82.975 248.015 83.295 ;
        RECT 248.215 82.975 248.475 83.295 ;
        RECT 246.895 81.595 247.035 82.895 ;
        RECT 247.295 82.295 247.555 82.615 ;
        RECT 246.835 81.275 247.095 81.595 ;
        RECT 246.375 80.595 246.635 80.915 ;
        RECT 243.615 80.430 243.875 80.575 ;
        RECT 243.605 80.060 243.885 80.430 ;
        RECT 244.075 80.255 244.335 80.575 ;
        RECT 244.535 79.915 244.795 80.235 ;
        RECT 244.595 79.750 244.735 79.915 ;
        RECT 244.525 79.380 244.805 79.750 ;
        RECT 245.455 79.575 245.715 79.895 ;
        RECT 246.375 79.575 246.635 79.895 ;
        RECT 244.075 77.875 244.335 78.195 ;
        RECT 244.135 77.710 244.275 77.875 ;
        RECT 244.065 77.340 244.345 77.710 ;
        RECT 243.615 75.835 243.875 76.155 ;
        RECT 243.675 74.795 243.815 75.835 ;
        RECT 243.615 74.475 243.875 74.795 ;
        RECT 243.155 73.115 243.415 73.435 ;
        RECT 243.215 71.590 243.355 73.115 ;
        RECT 243.675 72.755 243.815 74.475 ;
        RECT 243.615 72.435 243.875 72.755 ;
        RECT 243.145 71.220 243.425 71.590 ;
        RECT 243.675 70.230 243.815 72.435 ;
        RECT 243.605 69.860 243.885 70.230 ;
        RECT 244.135 67.995 244.275 77.340 ;
        RECT 244.595 70.035 244.735 79.380 ;
        RECT 245.515 78.535 245.655 79.575 ;
        RECT 245.455 78.215 245.715 78.535 ;
        RECT 246.435 77.855 246.575 79.575 ;
        RECT 247.355 78.195 247.495 82.295 ;
        RECT 247.815 81.595 247.955 82.975 ;
        RECT 247.755 81.275 248.015 81.595 ;
        RECT 248.275 80.430 248.415 82.975 ;
        RECT 249.195 82.470 249.335 85.695 ;
        RECT 250.505 85.500 250.785 85.870 ;
        RECT 250.055 85.015 250.315 85.335 ;
        RECT 249.125 82.100 249.405 82.470 ;
        RECT 249.595 82.295 249.855 82.615 ;
        RECT 248.675 81.275 248.935 81.595 ;
        RECT 248.205 80.060 248.485 80.430 ;
        RECT 247.755 79.575 248.015 79.895 ;
        RECT 247.295 77.875 247.555 78.195 ;
        RECT 246.375 77.535 246.635 77.855 ;
        RECT 247.815 75.135 247.955 79.575 ;
        RECT 248.735 78.535 248.875 81.275 ;
        RECT 249.655 80.575 249.795 82.295 ;
        RECT 249.595 80.255 249.855 80.575 ;
        RECT 248.675 78.215 248.935 78.535 ;
        RECT 248.215 76.855 248.475 77.175 ;
        RECT 248.275 75.815 248.415 76.855 ;
        RECT 248.215 75.495 248.475 75.815 ;
        RECT 244.995 74.815 245.255 75.135 ;
        RECT 247.755 74.815 248.015 75.135 ;
        RECT 244.535 69.715 244.795 70.035 ;
        RECT 244.535 69.035 244.795 69.355 ;
        RECT 244.075 67.675 244.335 67.995 ;
        RECT 242.755 67.085 243.815 67.225 ;
        RECT 242.295 66.575 242.895 66.715 ;
        RECT 241.775 65.975 242.035 66.295 ;
        RECT 242.235 65.975 242.495 66.295 ;
        RECT 242.295 65.275 242.435 65.975 ;
        RECT 241.315 64.955 241.575 65.275 ;
        RECT 242.235 64.955 242.495 65.275 ;
        RECT 242.235 62.235 242.495 62.555 ;
        RECT 239.925 58.980 240.205 59.350 ;
        RECT 242.295 59.155 242.435 62.235 ;
        RECT 242.235 58.835 242.495 59.155 ;
        RECT 242.755 58.475 242.895 66.575 ;
        RECT 243.155 63.935 243.415 64.255 ;
        RECT 243.215 62.555 243.355 63.935 ;
        RECT 243.675 62.555 243.815 67.085 ;
        RECT 244.595 66.975 244.735 69.035 ;
        RECT 244.535 66.655 244.795 66.975 ;
        RECT 244.525 65.780 244.805 66.150 ;
        RECT 244.075 64.615 244.335 64.935 ;
        RECT 244.135 63.430 244.275 64.615 ;
        RECT 244.595 64.255 244.735 65.780 ;
        RECT 244.535 63.935 244.795 64.255 ;
        RECT 244.065 63.060 244.345 63.430 ;
        RECT 243.155 62.235 243.415 62.555 ;
        RECT 243.615 62.235 243.875 62.555 ;
        RECT 243.675 61.875 243.815 62.235 ;
        RECT 244.135 61.875 244.275 63.060 ;
        RECT 243.615 61.555 243.875 61.875 ;
        RECT 244.075 61.555 244.335 61.875 ;
        RECT 244.535 61.555 244.795 61.875 ;
        RECT 242.695 58.155 242.955 58.475 ;
        RECT 243.675 58.135 243.815 61.555 ;
        RECT 239.475 57.815 239.735 58.135 ;
        RECT 243.615 57.815 243.875 58.135 ;
        RECT 239.015 56.115 239.275 56.435 ;
        RECT 239.075 45.215 239.215 56.115 ;
        RECT 239.535 51.335 239.675 57.815 ;
        RECT 242.235 56.115 242.495 56.435 ;
        RECT 239.935 55.095 240.195 55.415 ;
        RECT 241.775 55.095 242.035 55.415 ;
        RECT 239.475 51.015 239.735 51.335 ;
        RECT 239.995 48.275 240.135 55.095 ;
        RECT 241.835 53.375 241.975 55.095 ;
        RECT 241.775 53.055 242.035 53.375 ;
        RECT 241.315 52.375 241.575 52.695 ;
        RECT 241.375 50.995 241.515 52.375 ;
        RECT 241.315 50.675 241.575 50.995 ;
        RECT 241.375 48.615 241.515 50.675 ;
        RECT 242.295 48.955 242.435 56.115 ;
        RECT 243.155 55.435 243.415 55.755 ;
        RECT 242.695 52.715 242.955 53.035 ;
        RECT 242.755 50.995 242.895 52.715 ;
        RECT 243.215 50.995 243.355 55.435 ;
        RECT 244.595 53.910 244.735 61.555 ;
        RECT 244.525 53.540 244.805 53.910 ;
        RECT 245.055 53.795 245.195 74.815 ;
        RECT 250.115 73.095 250.255 85.015 ;
        RECT 250.575 83.635 250.715 85.500 ;
        RECT 250.515 83.315 250.775 83.635 ;
        RECT 250.575 79.895 250.715 83.315 ;
        RECT 252.415 81.110 252.555 86.375 ;
        RECT 253.335 86.265 253.475 108.815 ;
        RECT 253.795 105.735 253.935 109.225 ;
        RECT 254.655 108.135 254.915 108.455 ;
        RECT 253.735 105.415 253.995 105.735 ;
        RECT 254.715 102.335 254.855 108.135 ;
        RECT 255.115 104.055 255.375 104.375 ;
        RECT 255.175 102.675 255.315 104.055 ;
        RECT 255.115 102.355 255.375 102.675 ;
        RECT 254.185 101.820 254.465 102.190 ;
        RECT 254.655 102.015 254.915 102.335 ;
        RECT 254.255 96.895 254.395 101.820 ;
        RECT 254.715 97.575 254.855 102.015 ;
        RECT 256.095 100.715 256.235 109.225 ;
        RECT 258.395 107.435 258.535 109.225 ;
        RECT 259.715 108.475 259.975 108.795 ;
        RECT 257.875 107.115 258.135 107.435 ;
        RECT 258.335 107.115 258.595 107.435 ;
        RECT 257.935 105.395 258.075 107.115 ;
        RECT 259.775 105.395 259.915 108.475 ;
        RECT 257.875 105.075 258.135 105.395 ;
        RECT 259.715 105.075 259.975 105.395 ;
        RECT 257.415 104.055 257.675 104.375 ;
        RECT 257.475 103.355 257.615 104.055 ;
        RECT 257.415 103.035 257.675 103.355 ;
        RECT 257.415 102.015 257.675 102.335 ;
        RECT 257.935 102.190 258.075 105.075 ;
        RECT 258.795 104.735 259.055 105.055 ;
        RECT 260.175 104.735 260.435 105.055 ;
        RECT 258.855 104.375 258.995 104.735 ;
        RECT 258.795 104.055 259.055 104.375 ;
        RECT 256.095 100.575 256.695 100.715 ;
        RECT 257.475 100.635 257.615 102.015 ;
        RECT 257.865 101.820 258.145 102.190 ;
        RECT 260.235 101.995 260.375 104.735 ;
        RECT 260.695 103.355 260.835 109.225 ;
        RECT 261.555 107.795 261.815 108.115 ;
        RECT 261.615 105.395 261.755 107.795 ;
        RECT 262.015 107.455 262.275 107.775 ;
        RECT 262.075 105.395 262.215 107.455 ;
        RECT 261.555 105.075 261.815 105.395 ;
        RECT 262.015 105.075 262.275 105.395 ;
        RECT 260.635 103.035 260.895 103.355 ;
        RECT 260.175 101.675 260.435 101.995 ;
        RECT 257.875 101.335 258.135 101.655 ;
        RECT 256.555 99.275 256.695 100.575 ;
        RECT 257.415 100.315 257.675 100.635 ;
        RECT 257.935 100.295 258.075 101.335 ;
        RECT 257.875 99.975 258.135 100.295 ;
        RECT 256.955 99.295 257.215 99.615 ;
        RECT 256.495 98.955 256.755 99.275 ;
        RECT 257.015 97.915 257.155 99.295 ;
        RECT 257.405 98.420 257.685 98.790 ;
        RECT 258.335 98.615 258.595 98.935 ;
        RECT 256.955 97.595 257.215 97.915 ;
        RECT 254.655 97.255 254.915 97.575 ;
        RECT 257.475 96.895 257.615 98.420 ;
        RECT 258.395 96.895 258.535 98.615 ;
        RECT 260.235 97.575 260.375 101.675 ;
        RECT 262.075 99.615 262.215 105.075 ;
        RECT 262.475 99.635 262.735 99.955 ;
        RECT 262.015 99.295 262.275 99.615 ;
        RECT 260.175 97.255 260.435 97.575 ;
        RECT 253.735 96.575 253.995 96.895 ;
        RECT 254.195 96.575 254.455 96.895 ;
        RECT 257.415 96.635 257.675 96.895 ;
        RECT 257.415 96.575 258.075 96.635 ;
        RECT 258.335 96.575 258.595 96.895 ;
        RECT 258.795 96.575 259.055 96.895 ;
        RECT 253.795 91.795 253.935 96.575 ;
        RECT 254.655 96.235 254.915 96.555 ;
        RECT 257.475 96.495 258.075 96.575 ;
        RECT 254.715 94.175 254.855 96.235 ;
        RECT 257.935 96.215 258.075 96.495 ;
        RECT 255.105 95.700 255.385 96.070 ;
        RECT 257.875 95.895 258.135 96.215 ;
        RECT 255.175 94.855 255.315 95.700 ;
        RECT 255.115 94.535 255.375 94.855 ;
        RECT 254.655 93.855 254.915 94.175 ;
        RECT 253.735 91.475 253.995 91.795 ;
        RECT 254.715 89.835 254.855 93.855 ;
        RECT 255.175 90.630 255.315 94.535 ;
        RECT 257.875 93.855 258.135 94.175 ;
        RECT 257.935 91.795 258.075 93.855 ;
        RECT 257.875 91.475 258.135 91.795 ;
        RECT 257.415 91.135 257.675 91.455 ;
        RECT 255.105 90.260 255.385 90.630 ;
        RECT 252.875 86.125 253.475 86.265 ;
        RECT 253.795 89.695 254.855 89.835 ;
        RECT 252.345 80.740 252.625 81.110 ;
        RECT 252.875 80.575 253.015 86.125 ;
        RECT 253.275 85.355 253.535 85.675 ;
        RECT 253.335 83.975 253.475 85.355 ;
        RECT 253.275 83.655 253.535 83.975 ;
        RECT 252.815 80.255 253.075 80.575 ;
        RECT 250.515 79.575 250.775 79.895 ;
        RECT 253.795 73.395 253.935 89.695 ;
        RECT 255.175 89.325 255.315 90.260 ;
        RECT 254.715 89.185 255.315 89.325 ;
        RECT 254.195 80.255 254.455 80.575 ;
        RECT 252.875 73.255 253.935 73.395 ;
        RECT 250.055 72.775 250.315 73.095 ;
        RECT 245.915 72.435 246.175 72.755 ;
        RECT 246.835 72.435 247.095 72.755 ;
        RECT 245.975 72.270 246.115 72.435 ;
        RECT 245.905 71.900 246.185 72.270 ;
        RECT 245.455 69.375 245.715 69.695 ;
        RECT 245.515 59.495 245.655 69.375 ;
        RECT 245.975 66.150 246.115 71.900 ;
        RECT 246.365 69.180 246.645 69.550 ;
        RECT 246.375 69.035 246.635 69.180 ;
        RECT 245.905 65.780 246.185 66.150 ;
        RECT 246.375 65.975 246.635 66.295 ;
        RECT 246.435 61.535 246.575 65.975 ;
        RECT 246.895 65.275 247.035 72.435 ;
        RECT 252.875 72.415 253.015 73.255 ;
        RECT 252.815 72.095 253.075 72.415 ;
        RECT 253.275 72.095 253.535 72.415 ;
        RECT 249.135 71.755 249.395 72.075 ;
        RECT 248.205 70.540 248.485 70.910 ;
        RECT 247.285 69.860 247.565 70.230 ;
        RECT 246.835 64.955 247.095 65.275 ;
        RECT 247.355 64.255 247.495 69.860 ;
        RECT 248.275 69.695 248.415 70.540 ;
        RECT 248.665 69.860 248.945 70.230 ;
        RECT 248.735 69.695 248.875 69.860 ;
        RECT 249.195 69.695 249.335 71.755 ;
        RECT 253.335 70.910 253.475 72.095 ;
        RECT 253.795 71.735 253.935 73.255 ;
        RECT 253.735 71.415 253.995 71.735 ;
        RECT 253.265 70.540 253.545 70.910 ;
        RECT 248.215 69.375 248.475 69.695 ;
        RECT 248.675 69.375 248.935 69.695 ;
        RECT 249.135 69.375 249.395 69.695 ;
        RECT 253.335 67.995 253.475 70.540 ;
        RECT 253.795 69.355 253.935 71.415 ;
        RECT 253.735 69.035 253.995 69.355 ;
        RECT 254.255 69.015 254.395 80.255 ;
        RECT 254.715 72.075 254.855 89.185 ;
        RECT 256.495 86.035 256.755 86.355 ;
        RECT 255.115 85.355 255.375 85.675 ;
        RECT 255.175 81.255 255.315 85.355 ;
        RECT 255.565 81.420 255.845 81.790 ;
        RECT 255.115 80.935 255.375 81.255 ;
        RECT 255.175 80.575 255.315 80.935 ;
        RECT 255.635 80.575 255.775 81.420 ;
        RECT 256.555 80.915 256.695 86.035 ;
        RECT 257.475 83.975 257.615 91.135 ;
        RECT 257.935 86.435 258.075 91.475 ;
        RECT 258.395 89.415 258.535 96.575 ;
        RECT 258.855 95.390 258.995 96.575 ;
        RECT 258.785 95.020 259.065 95.390 ;
        RECT 262.015 92.155 262.275 92.475 ;
        RECT 259.705 90.940 259.985 91.310 ;
        RECT 261.095 91.195 261.355 91.455 ;
        RECT 260.695 91.135 261.355 91.195 ;
        RECT 259.775 90.775 259.915 90.940 ;
        RECT 260.175 90.795 260.435 91.115 ;
        RECT 260.695 91.055 261.295 91.135 ;
        RECT 259.715 90.455 259.975 90.775 ;
        RECT 258.335 89.095 258.595 89.415 ;
        RECT 259.715 89.095 259.975 89.415 ;
        RECT 258.395 87.035 258.535 89.095 ;
        RECT 259.255 88.590 259.515 88.735 ;
        RECT 259.245 88.475 259.525 88.590 ;
        RECT 258.855 88.335 259.525 88.475 ;
        RECT 258.335 86.715 258.595 87.035 ;
        RECT 257.935 86.295 258.535 86.435 ;
        RECT 257.415 83.655 257.675 83.975 ;
        RECT 256.955 83.315 257.215 83.635 ;
        RECT 257.015 81.595 257.155 83.315 ;
        RECT 256.955 81.275 257.215 81.595 ;
        RECT 257.475 81.255 257.615 83.655 ;
        RECT 256.495 80.595 256.755 80.915 ;
        RECT 256.945 80.740 257.225 81.110 ;
        RECT 257.415 80.935 257.675 81.255 ;
        RECT 255.115 80.255 255.375 80.575 ;
        RECT 255.575 80.315 255.835 80.575 ;
        RECT 255.575 80.255 256.235 80.315 ;
        RECT 255.635 80.175 256.235 80.255 ;
        RECT 256.555 80.235 256.695 80.595 ;
        RECT 257.015 80.575 257.155 80.740 ;
        RECT 256.955 80.255 257.215 80.575 ;
        RECT 257.875 80.255 258.135 80.575 ;
        RECT 254.655 71.755 254.915 72.075 ;
        RECT 256.095 70.035 256.235 80.175 ;
        RECT 256.495 79.915 256.755 80.235 ;
        RECT 256.555 78.535 256.695 79.915 ;
        RECT 256.495 78.215 256.755 78.535 ;
        RECT 256.495 77.195 256.755 77.515 ;
        RECT 256.555 72.755 256.695 77.195 ;
        RECT 257.935 74.795 258.075 80.255 ;
        RECT 258.395 77.175 258.535 86.295 ;
        RECT 258.335 76.855 258.595 77.175 ;
        RECT 258.335 75.835 258.595 76.155 ;
        RECT 257.875 74.475 258.135 74.795 ;
        RECT 258.395 74.195 258.535 75.835 ;
        RECT 258.855 75.135 258.995 88.335 ;
        RECT 259.245 88.220 259.525 88.335 ;
        RECT 259.775 88.055 259.915 89.095 ;
        RECT 259.715 87.735 259.975 88.055 ;
        RECT 259.775 82.955 259.915 87.735 ;
        RECT 259.715 82.635 259.975 82.955 ;
        RECT 260.235 80.915 260.375 90.795 ;
        RECT 260.695 86.355 260.835 91.055 ;
        RECT 261.095 90.455 261.355 90.775 ;
        RECT 261.155 89.755 261.295 90.455 ;
        RECT 261.095 89.435 261.355 89.755 ;
        RECT 261.555 89.435 261.815 89.755 ;
        RECT 260.635 86.035 260.895 86.355 ;
        RECT 261.095 83.315 261.355 83.635 ;
        RECT 260.635 82.295 260.895 82.615 ;
        RECT 260.175 80.595 260.435 80.915 ;
        RECT 259.255 80.255 259.515 80.575 ;
        RECT 258.795 74.815 259.055 75.135 ;
        RECT 257.935 74.055 258.535 74.195 ;
        RECT 257.935 72.755 258.075 74.055 ;
        RECT 258.855 73.005 258.995 74.815 ;
        RECT 259.315 74.455 259.455 80.255 ;
        RECT 260.695 78.875 260.835 82.295 ;
        RECT 261.155 81.255 261.295 83.315 ;
        RECT 261.095 80.935 261.355 81.255 ;
        RECT 261.085 79.380 261.365 79.750 ;
        RECT 260.635 78.555 260.895 78.875 ;
        RECT 260.635 77.535 260.895 77.855 ;
        RECT 259.715 76.855 259.975 77.175 ;
        RECT 259.255 74.135 259.515 74.455 ;
        RECT 259.775 74.310 259.915 76.855 ;
        RECT 259.705 73.940 259.985 74.310 ;
        RECT 259.255 73.005 259.515 73.095 ;
        RECT 258.855 72.865 259.515 73.005 ;
        RECT 259.255 72.775 259.515 72.865 ;
        RECT 256.495 72.435 256.755 72.755 ;
        RECT 257.875 72.435 258.135 72.755 ;
        RECT 258.335 72.435 258.595 72.755 ;
        RECT 258.395 72.270 258.535 72.435 ;
        RECT 258.325 71.900 258.605 72.270 ;
        RECT 258.335 71.755 258.595 71.900 ;
        RECT 256.035 69.715 256.295 70.035 ;
        RECT 259.775 69.695 259.915 73.940 ;
        RECT 260.695 72.755 260.835 77.535 ;
        RECT 261.155 75.475 261.295 79.380 ;
        RECT 261.095 75.155 261.355 75.475 ;
        RECT 261.615 75.135 261.755 89.435 ;
        RECT 262.075 88.055 262.215 92.155 ;
        RECT 262.015 87.735 262.275 88.055 ;
        RECT 262.015 82.635 262.275 82.955 ;
        RECT 262.075 78.875 262.215 82.635 ;
        RECT 262.535 80.575 262.675 99.635 ;
        RECT 262.995 97.575 263.135 109.225 ;
        RECT 263.395 109.155 263.655 109.475 ;
        RECT 265.225 109.225 265.505 132.985 ;
        RECT 267.525 109.225 267.805 133.565 ;
        RECT 269.825 109.225 270.105 134.145 ;
        RECT 272.125 109.225 272.405 134.725 ;
        RECT 274.425 109.225 274.705 135.305 ;
        RECT 276.725 109.225 277.005 135.885 ;
        RECT 277.255 109.415 278.315 109.555 ;
        RECT 262.935 97.255 263.195 97.575 ;
        RECT 262.925 88.900 263.205 89.270 ;
        RECT 262.935 88.755 263.195 88.900 ;
        RECT 263.455 83.295 263.595 109.155 ;
        RECT 264.315 106.775 264.575 107.095 ;
        RECT 264.375 104.375 264.515 106.775 ;
        RECT 264.775 105.075 265.035 105.395 ;
        RECT 264.315 104.055 264.575 104.375 ;
        RECT 263.855 99.635 264.115 99.955 ;
        RECT 263.915 95.195 264.055 99.635 ;
        RECT 264.315 99.295 264.575 99.615 ;
        RECT 264.375 97.915 264.515 99.295 ;
        RECT 264.315 97.595 264.575 97.915 ;
        RECT 263.855 94.875 264.115 95.195 ;
        RECT 263.915 88.395 264.055 94.875 ;
        RECT 264.835 91.195 264.975 105.075 ;
        RECT 265.295 97.915 265.435 109.225 ;
        RECT 266.155 104.735 266.415 105.055 ;
        RECT 266.215 103.015 266.355 104.735 ;
        RECT 267.595 104.715 267.735 109.225 ;
        RECT 269.895 106.155 270.035 109.225 ;
        RECT 272.195 107.775 272.335 109.225 ;
        RECT 272.135 107.455 272.395 107.775 ;
        RECT 269.895 106.015 270.495 106.155 ;
        RECT 270.355 105.735 270.495 106.015 ;
        RECT 270.295 105.415 270.555 105.735 ;
        RECT 268.455 105.075 268.715 105.395 ;
        RECT 270.755 105.075 271.015 105.395 ;
        RECT 267.535 104.395 267.795 104.715 ;
        RECT 266.155 102.695 266.415 103.015 ;
        RECT 265.235 97.595 265.495 97.915 ;
        RECT 265.235 93.855 265.495 94.175 ;
        RECT 265.295 91.455 265.435 93.855 ;
        RECT 266.215 92.475 266.355 102.695 ;
        RECT 267.995 101.675 268.255 101.995 ;
        RECT 268.055 100.635 268.195 101.675 ;
        RECT 267.995 100.315 268.255 100.635 ;
        RECT 266.155 92.155 266.415 92.475 ;
        RECT 266.215 91.795 266.355 92.155 ;
        RECT 266.155 91.475 266.415 91.795 ;
        RECT 264.375 91.055 264.975 91.195 ;
        RECT 265.235 91.135 265.495 91.455 ;
        RECT 267.535 91.135 267.795 91.455 ;
        RECT 263.855 88.075 264.115 88.395 ;
        RECT 264.375 83.715 264.515 91.055 ;
        RECT 266.615 90.795 266.875 91.115 ;
        RECT 267.075 90.795 267.335 91.115 ;
        RECT 264.775 90.455 265.035 90.775 ;
        RECT 264.835 84.395 264.975 90.455 ;
        RECT 265.235 88.985 265.495 89.075 ;
        RECT 265.235 88.845 266.355 88.985 ;
        RECT 265.235 88.755 265.495 88.845 ;
        RECT 264.835 84.255 265.895 84.395 ;
        RECT 264.375 83.575 264.975 83.715 ;
        RECT 263.395 82.975 263.655 83.295 ;
        RECT 262.935 82.295 263.195 82.615 ;
        RECT 262.475 80.255 262.735 80.575 ;
        RECT 262.015 78.555 262.275 78.875 ;
        RECT 262.015 77.875 262.275 78.195 ;
        RECT 262.075 77.175 262.215 77.875 ;
        RECT 262.015 76.855 262.275 77.175 ;
        RECT 261.555 74.815 261.815 75.135 ;
        RECT 261.095 74.135 261.355 74.455 ;
        RECT 260.635 72.435 260.895 72.755 ;
        RECT 260.165 71.220 260.445 71.590 ;
        RECT 260.235 70.715 260.375 71.220 ;
        RECT 260.175 70.395 260.435 70.715 ;
        RECT 257.415 69.375 257.675 69.695 ;
        RECT 259.255 69.375 259.515 69.695 ;
        RECT 259.715 69.375 259.975 69.695 ;
        RECT 254.195 68.695 254.455 69.015 ;
        RECT 253.275 67.675 253.535 67.995 ;
        RECT 248.215 67.335 248.475 67.655 ;
        RECT 247.295 63.935 247.555 64.255 ;
        RECT 248.275 62.555 248.415 67.335 ;
        RECT 248.675 66.655 248.935 66.975 ;
        RECT 248.215 62.235 248.475 62.555 ;
        RECT 247.755 61.895 248.015 62.215 ;
        RECT 248.735 61.955 248.875 66.655 ;
        RECT 252.345 63.740 252.625 64.110 ;
        RECT 256.955 63.935 257.215 64.255 ;
        RECT 252.415 62.555 252.555 63.740 ;
        RECT 252.355 62.235 252.615 62.555 ;
        RECT 255.575 62.235 255.835 62.555 ;
        RECT 246.835 61.555 247.095 61.875 ;
        RECT 246.375 61.215 246.635 61.535 ;
        RECT 246.435 60.855 246.575 61.215 ;
        RECT 246.375 60.535 246.635 60.855 ;
        RECT 245.455 59.175 245.715 59.495 ;
        RECT 246.435 58.815 246.575 60.535 ;
        RECT 246.375 58.495 246.635 58.815 ;
        RECT 245.915 58.155 246.175 58.475 ;
        RECT 245.975 53.910 246.115 58.155 ;
        RECT 246.435 54.055 246.575 58.495 ;
        RECT 246.895 54.590 247.035 61.555 ;
        RECT 247.815 56.435 247.955 61.895 ;
        RECT 248.275 61.815 248.875 61.955 ;
        RECT 248.275 60.855 248.415 61.815 ;
        RECT 252.815 61.555 253.075 61.875 ;
        RECT 248.215 60.535 248.475 60.855 ;
        RECT 248.275 59.155 248.415 60.535 ;
        RECT 252.875 59.835 253.015 61.555 ;
        RECT 255.635 60.855 255.775 62.235 ;
        RECT 257.015 61.195 257.155 63.935 ;
        RECT 257.475 61.955 257.615 69.375 ;
        RECT 259.315 69.015 259.455 69.375 ;
        RECT 259.255 68.695 259.515 69.015 ;
        RECT 257.875 66.655 258.135 66.975 ;
        RECT 257.935 62.555 258.075 66.655 ;
        RECT 257.875 62.235 258.135 62.555 ;
        RECT 257.475 61.815 258.075 61.955 ;
        RECT 257.415 61.390 257.675 61.535 ;
        RECT 256.955 60.875 257.215 61.195 ;
        RECT 257.405 61.020 257.685 61.390 ;
        RECT 254.655 60.535 254.915 60.855 ;
        RECT 255.115 60.535 255.375 60.855 ;
        RECT 255.575 60.535 255.835 60.855 ;
        RECT 252.815 59.515 253.075 59.835 ;
        RECT 248.215 58.835 248.475 59.155 ;
        RECT 254.195 58.835 254.455 59.155 ;
        RECT 248.275 58.135 248.415 58.835 ;
        RECT 248.215 57.815 248.475 58.135 ;
        RECT 248.215 56.455 248.475 56.775 ;
        RECT 252.815 56.455 253.075 56.775 ;
        RECT 247.755 56.115 248.015 56.435 ;
        RECT 248.275 55.835 248.415 56.455 ;
        RECT 252.355 56.115 252.615 56.435 ;
        RECT 247.355 55.695 248.415 55.835 ;
        RECT 250.975 55.775 251.235 56.095 ;
        RECT 246.825 54.220 247.105 54.590 ;
        RECT 245.055 53.655 245.655 53.795 ;
        RECT 244.995 53.055 245.255 53.375 ;
        RECT 244.535 52.715 244.795 53.035 ;
        RECT 242.695 50.675 242.955 50.995 ;
        RECT 243.155 50.675 243.415 50.995 ;
        RECT 242.235 48.635 242.495 48.955 ;
        RECT 241.315 48.295 241.575 48.615 ;
        RECT 239.935 47.955 240.195 48.275 ;
        RECT 241.375 45.555 241.515 48.295 ;
        RECT 242.295 45.895 242.435 48.635 ;
        RECT 242.235 45.575 242.495 45.895 ;
        RECT 242.755 45.555 242.895 50.675 ;
        RECT 244.595 49.035 244.735 52.715 ;
        RECT 245.055 49.975 245.195 53.055 ;
        RECT 244.995 49.655 245.255 49.975 ;
        RECT 244.595 48.895 245.195 49.035 ;
        RECT 243.155 47.615 243.415 47.935 ;
        RECT 243.215 46.235 243.355 47.615 ;
        RECT 245.055 47.255 245.195 48.895 ;
        RECT 244.995 46.935 245.255 47.255 ;
        RECT 243.155 45.915 243.415 46.235 ;
        RECT 241.315 45.235 241.575 45.555 ;
        RECT 242.695 45.235 242.955 45.555 ;
        RECT 239.015 44.895 239.275 45.215 ;
        RECT 238.555 41.495 238.815 41.815 ;
        RECT 237.175 40.475 237.435 40.795 ;
        RECT 238.615 40.115 238.755 41.495 ;
        RECT 238.555 39.795 238.815 40.115 ;
        RECT 239.075 39.775 239.215 44.895 ;
        RECT 242.755 43.595 242.895 45.235 ;
        RECT 242.295 43.455 242.895 43.595 ;
        RECT 242.295 42.835 242.435 43.455 ;
        RECT 242.695 42.855 242.955 43.175 ;
        RECT 242.235 42.515 242.495 42.835 ;
        RECT 242.235 41.495 242.495 41.815 ;
        RECT 242.295 40.795 242.435 41.495 ;
        RECT 242.235 40.475 242.495 40.795 ;
        RECT 239.015 39.455 239.275 39.775 ;
        RECT 241.315 38.775 241.575 39.095 ;
        RECT 242.235 38.775 242.495 39.095 ;
        RECT 241.375 36.715 241.515 38.775 ;
        RECT 236.715 36.395 236.975 36.715 ;
        RECT 241.315 36.395 241.575 36.715 ;
        RECT 236.775 35.355 236.915 36.395 ;
        RECT 233.495 35.035 233.755 35.355 ;
        RECT 236.715 35.035 236.975 35.355 ;
        RECT 242.295 35.015 242.435 38.775 ;
        RECT 242.235 34.695 242.495 35.015 ;
        RECT 232.575 34.355 232.835 34.675 ;
        RECT 242.235 34.015 242.495 34.335 ;
        RECT 242.295 32.635 242.435 34.015 ;
        RECT 242.755 32.635 242.895 42.855 ;
        RECT 243.215 42.235 243.355 45.915 ;
        RECT 244.535 44.555 244.795 44.875 ;
        RECT 244.595 42.835 244.735 44.555 ;
        RECT 244.535 42.515 244.795 42.835 ;
        RECT 245.055 42.495 245.195 46.935 ;
        RECT 243.215 42.095 243.815 42.235 ;
        RECT 244.995 42.175 245.255 42.495 ;
        RECT 243.155 41.495 243.415 41.815 ;
        RECT 242.235 32.315 242.495 32.635 ;
        RECT 242.695 32.315 242.955 32.635 ;
        RECT 216.475 31.295 216.735 31.615 ;
        RECT 219.235 31.295 219.495 31.615 ;
        RECT 227.975 31.295 228.235 31.615 ;
        RECT 243.215 30.935 243.355 41.495 ;
        RECT 243.675 38.835 243.815 42.095 ;
        RECT 245.515 40.455 245.655 53.655 ;
        RECT 245.905 53.540 246.185 53.910 ;
        RECT 246.375 53.735 246.635 54.055 ;
        RECT 246.375 51.015 246.635 51.335 ;
        RECT 246.435 50.655 246.575 51.015 ;
        RECT 247.355 50.995 247.495 55.695 ;
        RECT 249.135 52.375 249.395 52.695 ;
        RECT 249.195 50.995 249.335 52.375 ;
        RECT 247.295 50.675 247.555 50.995 ;
        RECT 247.755 50.675 248.015 50.995 ;
        RECT 249.135 50.675 249.395 50.995 ;
        RECT 246.375 50.335 246.635 50.655 ;
        RECT 247.815 48.955 247.955 50.675 ;
        RECT 249.595 49.655 249.855 49.975 ;
        RECT 247.755 48.635 248.015 48.955 ;
        RECT 248.675 47.275 248.935 47.595 ;
        RECT 246.375 45.235 246.635 45.555 ;
        RECT 246.435 43.175 246.575 45.235 ;
        RECT 248.735 43.515 248.875 47.275 ;
        RECT 249.655 45.215 249.795 49.655 ;
        RECT 250.055 47.615 250.315 47.935 ;
        RECT 250.115 45.895 250.255 47.615 ;
        RECT 250.055 45.575 250.315 45.895 ;
        RECT 249.595 44.895 249.855 45.215 ;
        RECT 248.675 43.195 248.935 43.515 ;
        RECT 245.915 42.855 246.175 43.175 ;
        RECT 246.375 42.855 246.635 43.175 ;
        RECT 245.455 40.135 245.715 40.455 ;
        RECT 243.675 38.695 244.275 38.835 ;
        RECT 244.135 36.715 244.275 38.695 ;
        RECT 244.535 37.075 244.795 37.395 ;
        RECT 244.075 36.395 244.335 36.715 ;
        RECT 244.135 35.015 244.275 36.395 ;
        RECT 244.075 34.755 244.335 35.015 ;
        RECT 243.675 34.695 244.335 34.755 ;
        RECT 243.675 34.615 244.275 34.695 ;
        RECT 243.675 31.275 243.815 34.615 ;
        RECT 244.595 33.655 244.735 37.075 ;
        RECT 245.515 36.375 245.655 40.135 ;
        RECT 245.975 39.095 246.115 42.855 ;
        RECT 251.035 42.495 251.175 55.775 ;
        RECT 252.415 54.395 252.555 56.115 ;
        RECT 252.355 54.075 252.615 54.395 ;
        RECT 252.875 53.715 253.015 56.455 ;
        RECT 254.255 56.095 254.395 58.835 ;
        RECT 254.715 58.475 254.855 60.535 ;
        RECT 254.655 58.155 254.915 58.475 ;
        RECT 255.175 56.775 255.315 60.535 ;
        RECT 257.935 59.155 258.075 61.815 ;
        RECT 259.315 59.835 259.455 68.695 ;
        RECT 259.775 67.315 259.915 69.375 ;
        RECT 260.695 68.925 260.835 72.435 ;
        RECT 261.155 69.695 261.295 74.135 ;
        RECT 261.615 70.035 261.755 74.815 ;
        RECT 262.075 70.035 262.215 76.855 ;
        RECT 262.535 76.350 262.675 80.255 ;
        RECT 262.465 75.980 262.745 76.350 ;
        RECT 262.475 75.495 262.735 75.815 ;
        RECT 261.555 69.715 261.815 70.035 ;
        RECT 262.015 69.715 262.275 70.035 ;
        RECT 261.095 69.375 261.355 69.695 ;
        RECT 262.015 69.035 262.275 69.355 ;
        RECT 260.695 68.785 261.295 68.925 ;
        RECT 259.715 66.995 259.975 67.315 ;
        RECT 259.775 65.275 259.915 66.995 ;
        RECT 259.715 64.955 259.975 65.275 ;
        RECT 260.175 64.955 260.435 65.275 ;
        RECT 259.775 61.875 259.915 64.955 ;
        RECT 260.235 62.750 260.375 64.955 ;
        RECT 260.625 64.420 260.905 64.790 ;
        RECT 260.695 63.915 260.835 64.420 ;
        RECT 260.635 63.595 260.895 63.915 ;
        RECT 260.165 62.380 260.445 62.750 ;
        RECT 260.695 62.555 260.835 63.595 ;
        RECT 259.715 61.555 259.975 61.875 ;
        RECT 260.235 60.855 260.375 62.380 ;
        RECT 260.635 62.235 260.895 62.555 ;
        RECT 260.175 60.535 260.435 60.855 ;
        RECT 259.255 59.515 259.515 59.835 ;
        RECT 257.875 58.835 258.135 59.155 ;
        RECT 258.325 58.980 258.605 59.350 ;
        RECT 255.115 56.455 255.375 56.775 ;
        RECT 254.195 55.775 254.455 56.095 ;
        RECT 257.875 55.775 258.135 56.095 ;
        RECT 252.815 53.395 253.075 53.715 ;
        RECT 254.255 53.035 254.395 55.775 ;
        RECT 257.415 55.095 257.675 55.415 ;
        RECT 254.195 52.715 254.455 53.035 ;
        RECT 255.575 52.715 255.835 53.035 ;
        RECT 255.635 50.655 255.775 52.715 ;
        RECT 257.475 51.335 257.615 55.095 ;
        RECT 257.935 52.695 258.075 55.775 ;
        RECT 258.395 53.375 258.535 58.980 ;
        RECT 260.635 58.155 260.895 58.475 ;
        RECT 260.695 56.775 260.835 58.155 ;
        RECT 260.635 56.455 260.895 56.775 ;
        RECT 258.335 53.055 258.595 53.375 ;
        RECT 258.795 52.715 259.055 53.035 ;
        RECT 257.875 52.375 258.135 52.695 ;
        RECT 256.035 51.015 256.295 51.335 ;
        RECT 257.415 51.015 257.675 51.335 ;
        RECT 255.575 50.335 255.835 50.655 ;
        RECT 254.655 48.635 254.915 48.955 ;
        RECT 251.895 46.935 252.155 47.255 ;
        RECT 251.955 45.895 252.095 46.935 ;
        RECT 251.895 45.575 252.155 45.895 ;
        RECT 254.715 45.215 254.855 48.635 ;
        RECT 255.635 47.935 255.775 50.335 ;
        RECT 255.575 47.615 255.835 47.935 ;
        RECT 255.575 46.935 255.835 47.255 ;
        RECT 254.655 44.895 254.915 45.215 ;
        RECT 250.975 42.175 251.235 42.495 ;
        RECT 254.715 40.455 254.855 44.895 ;
        RECT 255.635 44.535 255.775 46.935 ;
        RECT 255.575 44.215 255.835 44.535 ;
        RECT 256.095 43.515 256.235 51.015 ;
        RECT 257.415 47.275 257.675 47.595 ;
        RECT 257.475 46.235 257.615 47.275 ;
        RECT 257.415 45.915 257.675 46.235 ;
        RECT 256.955 44.555 257.215 44.875 ;
        RECT 256.035 43.195 256.295 43.515 ;
        RECT 256.035 42.175 256.295 42.495 ;
        RECT 254.655 40.135 254.915 40.455 ;
        RECT 252.355 39.455 252.615 39.775 ;
        RECT 245.915 38.775 246.175 39.095 ;
        RECT 245.455 36.055 245.715 36.375 ;
        RECT 245.975 34.755 246.115 38.775 ;
        RECT 252.415 35.355 252.555 39.455 ;
        RECT 256.095 37.395 256.235 42.175 ;
        RECT 257.015 42.155 257.155 44.555 ;
        RECT 258.855 42.495 258.995 52.715 ;
        RECT 260.695 51.675 260.835 56.455 ;
        RECT 261.155 55.155 261.295 68.785 ;
        RECT 262.075 67.995 262.215 69.035 ;
        RECT 262.015 67.675 262.275 67.995 ;
        RECT 262.535 66.975 262.675 75.495 ;
        RECT 262.995 71.590 263.135 82.295 ;
        RECT 263.455 75.815 263.595 82.975 ;
        RECT 263.855 80.255 264.115 80.575 ;
        RECT 263.395 75.495 263.655 75.815 ;
        RECT 263.385 74.620 263.665 74.990 ;
        RECT 263.455 73.095 263.595 74.620 ;
        RECT 263.395 72.775 263.655 73.095 ;
        RECT 262.925 71.220 263.205 71.590 ;
        RECT 263.915 70.115 264.055 80.255 ;
        RECT 264.315 77.535 264.575 77.855 ;
        RECT 264.375 76.155 264.515 77.535 ;
        RECT 264.315 75.835 264.575 76.155 ;
        RECT 264.315 74.815 264.575 75.135 ;
        RECT 264.375 72.755 264.515 74.815 ;
        RECT 264.835 72.950 264.975 83.575 ;
        RECT 265.235 83.315 265.495 83.635 ;
        RECT 265.295 78.535 265.435 83.315 ;
        RECT 265.235 78.215 265.495 78.535 ;
        RECT 265.755 73.395 265.895 84.255 ;
        RECT 266.215 81.255 266.355 88.845 ;
        RECT 266.675 85.675 266.815 90.795 ;
        RECT 267.135 89.075 267.275 90.795 ;
        RECT 267.075 88.755 267.335 89.075 ;
        RECT 267.135 88.395 267.275 88.755 ;
        RECT 267.075 88.075 267.335 88.395 ;
        RECT 267.595 86.695 267.735 91.135 ;
        RECT 267.535 86.375 267.795 86.695 ;
        RECT 266.615 85.355 266.875 85.675 ;
        RECT 266.675 83.635 266.815 85.355 ;
        RECT 266.615 83.315 266.875 83.635 ;
        RECT 266.155 81.110 266.415 81.255 ;
        RECT 266.145 80.740 266.425 81.110 ;
        RECT 267.595 80.995 267.735 86.375 ;
        RECT 268.515 81.505 268.655 105.075 ;
        RECT 268.915 104.395 269.175 104.715 ;
        RECT 268.975 100.635 269.115 104.395 ;
        RECT 269.835 102.355 270.095 102.675 ;
        RECT 268.915 100.315 269.175 100.635 ;
        RECT 269.365 100.460 269.645 100.830 ;
        RECT 269.435 99.615 269.575 100.460 ;
        RECT 269.375 99.295 269.635 99.615 ;
        RECT 269.895 99.525 270.035 102.355 ;
        RECT 270.295 99.525 270.555 99.615 ;
        RECT 269.895 99.385 270.555 99.525 ;
        RECT 268.915 90.455 269.175 90.775 ;
        RECT 268.975 89.075 269.115 90.455 ;
        RECT 268.915 88.755 269.175 89.075 ;
        RECT 269.895 86.355 270.035 99.385 ;
        RECT 270.295 99.295 270.555 99.385 ;
        RECT 270.815 88.475 270.955 105.075 ;
        RECT 274.495 101.995 274.635 109.225 ;
        RECT 276.795 108.875 276.935 109.225 ;
        RECT 277.255 108.875 277.395 109.415 ;
        RECT 276.795 108.735 277.395 108.875 ;
        RECT 276.735 107.115 276.995 107.435 ;
        RECT 276.795 106.075 276.935 107.115 ;
        RECT 276.735 105.755 276.995 106.075 ;
        RECT 275.355 104.735 275.615 105.055 ;
        RECT 274.435 101.675 274.695 101.995 ;
        RECT 275.415 101.655 275.555 104.735 ;
        RECT 277.195 104.055 277.455 104.375 ;
        RECT 277.255 102.335 277.395 104.055 ;
        RECT 277.195 102.015 277.455 102.335 ;
        RECT 275.355 101.335 275.615 101.655 ;
        RECT 273.055 99.295 273.315 99.615 ;
        RECT 273.115 97.915 273.255 99.295 ;
        RECT 273.055 97.595 273.315 97.915 ;
        RECT 275.415 97.235 275.555 101.335 ;
        RECT 276.735 98.615 276.995 98.935 ;
        RECT 276.795 97.235 276.935 98.615 ;
        RECT 275.355 96.915 275.615 97.235 ;
        RECT 276.735 96.915 276.995 97.235 ;
        RECT 277.255 96.895 277.395 102.015 ;
        RECT 277.655 101.335 277.915 101.655 ;
        RECT 277.715 100.635 277.855 101.335 ;
        RECT 277.655 100.315 277.915 100.635 ;
        RECT 272.595 96.575 272.855 96.895 ;
        RECT 276.275 96.750 276.535 96.895 ;
        RECT 271.215 89.095 271.475 89.415 ;
        RECT 270.355 88.335 270.955 88.475 ;
        RECT 269.835 86.035 270.095 86.355 ;
        RECT 269.895 83.635 270.035 86.035 ;
        RECT 270.355 85.335 270.495 88.335 ;
        RECT 270.755 87.735 271.015 88.055 ;
        RECT 270.295 85.015 270.555 85.335 ;
        RECT 269.835 83.315 270.095 83.635 ;
        RECT 269.375 82.295 269.635 82.615 ;
        RECT 267.135 80.855 267.735 80.995 ;
        RECT 268.055 81.365 268.655 81.505 ;
        RECT 267.135 80.575 267.275 80.855 ;
        RECT 266.155 80.430 266.415 80.575 ;
        RECT 266.145 80.060 266.425 80.430 ;
        RECT 267.075 80.255 267.335 80.575 ;
        RECT 267.535 80.255 267.795 80.575 ;
        RECT 266.615 74.135 266.875 74.455 ;
        RECT 265.755 73.255 266.355 73.395 ;
        RECT 264.315 72.435 264.575 72.755 ;
        RECT 264.765 72.580 265.045 72.950 ;
        RECT 265.695 72.775 265.955 73.095 ;
        RECT 265.235 72.435 265.495 72.755 ;
        RECT 265.295 72.155 265.435 72.435 ;
        RECT 265.755 72.270 265.895 72.775 ;
        RECT 262.995 69.975 264.055 70.115 ;
        RECT 264.835 72.015 265.435 72.155 ;
        RECT 262.475 66.655 262.735 66.975 ;
        RECT 262.535 55.755 262.675 66.655 ;
        RECT 262.995 58.815 263.135 69.975 ;
        RECT 264.315 69.715 264.575 70.035 ;
        RECT 263.855 69.375 264.115 69.695 ;
        RECT 264.375 69.550 264.515 69.715 ;
        RECT 263.915 67.655 264.055 69.375 ;
        RECT 264.305 69.180 264.585 69.550 ;
        RECT 263.855 67.335 264.115 67.655 ;
        RECT 264.835 66.635 264.975 72.015 ;
        RECT 265.685 71.900 265.965 72.270 ;
        RECT 265.695 71.415 265.955 71.735 ;
        RECT 265.755 70.715 265.895 71.415 ;
        RECT 265.695 70.395 265.955 70.715 ;
        RECT 266.215 67.995 266.355 73.255 ;
        RECT 266.675 69.695 266.815 74.135 ;
        RECT 267.595 73.395 267.735 80.255 ;
        RECT 268.055 78.195 268.195 81.365 ;
        RECT 268.455 80.595 268.715 80.915 ;
        RECT 268.515 78.875 268.655 80.595 ;
        RECT 269.435 80.575 269.575 82.295 ;
        RECT 270.355 81.595 270.495 85.015 ;
        RECT 270.295 81.275 270.555 81.595 ;
        RECT 269.375 80.255 269.635 80.575 ;
        RECT 268.915 79.915 269.175 80.235 ;
        RECT 268.455 78.555 268.715 78.875 ;
        RECT 267.995 77.875 268.255 78.195 ;
        RECT 268.055 74.795 268.195 77.875 ;
        RECT 268.975 77.595 269.115 79.915 ;
        RECT 270.295 79.575 270.555 79.895 ;
        RECT 270.355 78.390 270.495 79.575 ;
        RECT 270.285 78.020 270.565 78.390 ;
        RECT 268.515 77.515 269.115 77.595 ;
        RECT 268.455 77.455 269.115 77.515 ;
        RECT 268.455 77.195 268.715 77.455 ;
        RECT 267.995 74.475 268.255 74.795 ;
        RECT 267.595 73.255 268.195 73.395 ;
        RECT 268.055 72.755 268.195 73.255 ;
        RECT 268.975 72.755 269.115 77.455 ;
        RECT 270.815 73.435 270.955 87.735 ;
        RECT 270.755 73.115 271.015 73.435 ;
        RECT 267.995 72.435 268.255 72.755 ;
        RECT 268.915 72.435 269.175 72.755 ;
        RECT 267.535 71.755 267.795 72.075 ;
        RECT 267.595 70.715 267.735 71.755 ;
        RECT 268.055 70.715 268.195 72.435 ;
        RECT 268.455 71.755 268.715 72.075 ;
        RECT 267.535 70.395 267.795 70.715 ;
        RECT 267.995 70.395 268.255 70.715 ;
        RECT 268.515 69.695 268.655 71.755 ;
        RECT 266.615 69.375 266.875 69.695 ;
        RECT 268.455 69.375 268.715 69.695 ;
        RECT 266.615 68.695 266.875 69.015 ;
        RECT 269.375 68.695 269.635 69.015 ;
        RECT 266.675 68.190 266.815 68.695 ;
        RECT 266.155 67.675 266.415 67.995 ;
        RECT 266.605 67.820 266.885 68.190 ;
        RECT 269.435 67.510 269.575 68.695 ;
        RECT 269.365 67.140 269.645 67.510 ;
        RECT 271.275 66.635 271.415 89.095 ;
        RECT 272.655 77.855 272.795 96.575 ;
        RECT 276.265 96.380 276.545 96.750 ;
        RECT 277.195 96.635 277.455 96.895 ;
        RECT 276.795 96.575 277.455 96.635 ;
        RECT 276.795 96.495 277.395 96.575 ;
        RECT 275.815 95.955 276.075 96.215 ;
        RECT 273.575 95.895 276.075 95.955 ;
        RECT 273.575 95.815 276.015 95.895 ;
        RECT 273.575 93.835 273.715 95.815 ;
        RECT 276.795 94.515 276.935 96.495 ;
        RECT 277.185 95.020 277.465 95.390 ;
        RECT 277.715 95.195 277.855 100.315 ;
        RECT 278.175 99.355 278.315 109.415 ;
        RECT 279.025 109.225 279.305 136.465 ;
        RECT 281.325 109.225 281.605 137.045 ;
        RECT 283.625 109.225 283.905 137.625 ;
        RECT 285.925 109.225 286.205 138.205 ;
        RECT 288.225 109.225 288.505 138.785 ;
        RECT 290.525 109.225 290.805 139.365 ;
        RECT 292.825 109.225 293.105 139.945 ;
        RECT 295.125 109.225 295.405 140.525 ;
        RECT 295.655 109.415 297.175 109.555 ;
        RECT 279.095 107.095 279.235 109.225 ;
        RECT 279.035 106.775 279.295 107.095 ;
        RECT 279.035 105.075 279.295 105.395 ;
        RECT 280.415 105.075 280.675 105.395 ;
        RECT 278.175 99.275 278.775 99.355 ;
        RECT 278.175 99.215 278.835 99.275 ;
        RECT 278.575 98.955 278.835 99.215 ;
        RECT 279.095 98.935 279.235 105.075 ;
        RECT 280.475 102.335 280.615 105.075 ;
        RECT 280.415 102.015 280.675 102.335 ;
        RECT 280.475 100.295 280.615 102.015 ;
        RECT 280.865 101.820 281.145 102.190 ;
        RECT 280.415 99.975 280.675 100.295 ;
        RECT 280.935 99.955 281.075 101.820 ;
        RECT 281.395 100.295 281.535 109.225 ;
        RECT 282.715 107.455 282.975 107.775 ;
        RECT 282.255 104.735 282.515 105.055 ;
        RECT 281.795 100.315 282.055 100.635 ;
        RECT 281.335 99.975 281.595 100.295 ;
        RECT 280.875 99.635 281.135 99.955 ;
        RECT 279.035 98.615 279.295 98.935 ;
        RECT 278.575 96.235 278.835 96.555 ;
        RECT 277.255 94.515 277.395 95.020 ;
        RECT 277.655 94.875 277.915 95.195 ;
        RECT 278.635 94.515 278.775 96.235 ;
        RECT 279.095 96.215 279.235 98.615 ;
        RECT 279.945 97.740 280.225 98.110 ;
        RECT 280.015 97.235 280.155 97.740 ;
        RECT 279.495 96.915 279.755 97.235 ;
        RECT 279.955 96.915 280.215 97.235 ;
        RECT 279.035 95.895 279.295 96.215 ;
        RECT 279.555 95.195 279.695 96.915 ;
        RECT 280.015 96.215 280.155 96.915 ;
        RECT 279.955 95.895 280.215 96.215 ;
        RECT 279.495 94.875 279.755 95.195 ;
        RECT 280.875 94.535 281.135 94.855 ;
        RECT 276.735 94.195 276.995 94.515 ;
        RECT 277.195 94.195 277.455 94.515 ;
        RECT 278.575 94.195 278.835 94.515 ;
        RECT 273.515 93.515 273.775 93.835 ;
        RECT 274.435 93.175 274.695 93.495 ;
        RECT 274.495 89.415 274.635 93.175 ;
        RECT 279.955 92.155 280.215 92.475 ;
        RECT 280.015 91.455 280.155 92.155 ;
        RECT 280.935 91.455 281.075 94.535 ;
        RECT 281.855 91.795 281.995 100.315 ;
        RECT 282.315 97.915 282.455 104.735 ;
        RECT 282.775 98.935 282.915 107.455 ;
        RECT 282.715 98.615 282.975 98.935 ;
        RECT 283.695 97.915 283.835 109.225 ;
        RECT 285.995 102.755 286.135 109.225 ;
        RECT 285.995 102.615 287.055 102.755 ;
        RECT 285.935 101.675 286.195 101.995 ;
        RECT 285.995 100.635 286.135 101.675 ;
        RECT 285.935 100.315 286.195 100.635 ;
        RECT 285.475 99.635 285.735 99.955 ;
        RECT 286.395 99.635 286.655 99.955 ;
        RECT 282.255 97.595 282.515 97.915 ;
        RECT 283.635 97.595 283.895 97.915 ;
        RECT 283.635 96.915 283.895 97.235 ;
        RECT 282.715 96.575 282.975 96.895 ;
        RECT 282.775 94.515 282.915 96.575 ;
        RECT 283.175 96.235 283.435 96.555 ;
        RECT 283.235 94.515 283.375 96.235 ;
        RECT 282.715 94.195 282.975 94.515 ;
        RECT 283.175 94.195 283.435 94.515 ;
        RECT 281.795 91.475 282.055 91.795 ;
        RECT 278.115 91.135 278.375 91.455 ;
        RECT 279.955 91.135 280.215 91.455 ;
        RECT 280.875 91.135 281.135 91.455 ;
        RECT 274.435 89.095 274.695 89.415 ;
        RECT 276.275 86.715 276.535 87.035 ;
        RECT 276.335 83.975 276.475 86.715 ;
        RECT 276.275 83.655 276.535 83.975 ;
        RECT 274.435 82.975 274.695 83.295 ;
        RECT 272.595 77.535 272.855 77.855 ;
        RECT 272.135 72.775 272.395 73.095 ;
        RECT 272.195 71.735 272.335 72.775 ;
        RECT 272.135 71.415 272.395 71.735 ;
        RECT 272.195 70.035 272.335 71.415 ;
        RECT 272.135 69.715 272.395 70.035 ;
        RECT 274.495 69.695 274.635 82.975 ;
        RECT 276.335 81.505 276.475 83.655 ;
        RECT 278.175 83.635 278.315 91.135 ;
        RECT 279.035 90.795 279.295 91.115 ;
        RECT 278.575 90.455 278.835 90.775 ;
        RECT 278.635 88.055 278.775 90.455 ;
        RECT 279.095 89.075 279.235 90.795 ;
        RECT 279.495 90.455 279.755 90.775 ;
        RECT 279.035 88.755 279.295 89.075 ;
        RECT 278.575 87.735 278.835 88.055 ;
        RECT 278.115 83.545 278.375 83.635 ;
        RECT 275.875 81.365 276.475 81.505 ;
        RECT 277.715 83.405 278.375 83.545 ;
        RECT 275.875 75.135 276.015 81.365 ;
        RECT 276.275 75.155 276.535 75.475 ;
        RECT 275.815 74.815 276.075 75.135 ;
        RECT 276.335 72.415 276.475 75.155 ;
        RECT 277.195 74.705 277.455 74.795 ;
        RECT 277.715 74.705 277.855 83.405 ;
        RECT 278.115 83.315 278.375 83.405 ;
        RECT 277.195 74.565 277.855 74.705 ;
        RECT 277.195 74.475 277.455 74.565 ;
        RECT 276.275 72.095 276.535 72.415 ;
        RECT 272.595 69.375 272.855 69.695 ;
        RECT 274.435 69.375 274.695 69.695 ;
        RECT 272.655 67.315 272.795 69.375 ;
        RECT 273.055 69.035 273.315 69.355 ;
        RECT 273.115 67.315 273.255 69.035 ;
        RECT 272.595 66.995 272.855 67.315 ;
        RECT 273.055 66.995 273.315 67.315 ;
        RECT 264.775 66.315 265.035 66.635 ;
        RECT 271.215 66.315 271.475 66.635 ;
        RECT 263.395 64.615 263.655 64.935 ;
        RECT 263.455 58.815 263.595 64.615 ;
        RECT 271.275 63.575 271.415 66.315 ;
        RECT 272.655 63.915 272.795 66.995 ;
        RECT 273.115 65.275 273.255 66.995 ;
        RECT 273.055 64.955 273.315 65.275 ;
        RECT 274.495 63.915 274.635 69.375 ;
        RECT 276.335 66.295 276.475 72.095 ;
        RECT 277.715 67.655 277.855 74.565 ;
        RECT 278.115 74.475 278.375 74.795 ;
        RECT 279.025 74.620 279.305 74.990 ;
        RECT 278.175 72.755 278.315 74.475 ;
        RECT 279.095 74.455 279.235 74.620 ;
        RECT 279.035 74.135 279.295 74.455 ;
        RECT 278.115 72.435 278.375 72.755 ;
        RECT 277.655 67.335 277.915 67.655 ;
        RECT 278.175 66.975 278.315 72.435 ;
        RECT 278.575 72.095 278.835 72.415 ;
        RECT 278.635 69.695 278.775 72.095 ;
        RECT 278.575 69.375 278.835 69.695 ;
        RECT 278.115 66.655 278.375 66.975 ;
        RECT 276.275 65.975 276.535 66.295 ;
        RECT 276.335 64.255 276.475 65.975 ;
        RECT 278.175 64.595 278.315 66.655 ;
        RECT 278.635 64.595 278.775 69.375 ;
        RECT 279.555 64.935 279.695 90.455 ;
        RECT 280.415 87.735 280.675 88.055 ;
        RECT 280.475 83.830 280.615 87.735 ;
        RECT 283.695 86.355 283.835 96.915 ;
        RECT 284.555 96.575 284.815 96.895 ;
        RECT 283.635 86.265 283.895 86.355 ;
        RECT 282.775 86.125 283.895 86.265 ;
        RECT 280.405 83.460 280.685 83.830 ;
        RECT 279.955 80.935 280.215 81.255 ;
        RECT 280.015 73.095 280.155 80.935 ;
        RECT 280.415 80.255 280.675 80.575 ;
        RECT 280.475 78.875 280.615 80.255 ;
        RECT 281.335 79.575 281.595 79.895 ;
        RECT 280.415 78.555 280.675 78.875 ;
        RECT 281.395 73.395 281.535 79.575 ;
        RECT 280.935 73.255 281.535 73.395 ;
        RECT 279.955 72.775 280.215 73.095 ;
        RECT 279.955 69.035 280.215 69.355 ;
        RECT 280.015 67.995 280.155 69.035 ;
        RECT 279.955 67.675 280.215 67.995 ;
        RECT 280.415 67.675 280.675 67.995 ;
        RECT 280.475 66.830 280.615 67.675 ;
        RECT 280.405 66.460 280.685 66.830 ;
        RECT 279.495 64.615 279.755 64.935 ;
        RECT 278.115 64.275 278.375 64.595 ;
        RECT 278.575 64.275 278.835 64.595 ;
        RECT 276.275 63.935 276.535 64.255 ;
        RECT 272.595 63.595 272.855 63.915 ;
        RECT 274.435 63.595 274.695 63.915 ;
        RECT 270.755 63.255 271.015 63.575 ;
        RECT 271.215 63.255 271.475 63.575 ;
        RECT 270.815 62.555 270.955 63.255 ;
        RECT 270.755 62.235 271.015 62.555 ;
        RECT 274.495 62.215 274.635 63.595 ;
        RECT 274.435 61.895 274.695 62.215 ;
        RECT 274.495 58.815 274.635 61.895 ;
        RECT 276.335 61.875 276.475 63.935 ;
        RECT 278.175 62.215 278.315 64.275 ;
        RECT 280.935 62.555 281.075 73.255 ;
        RECT 282.245 72.580 282.525 72.950 ;
        RECT 281.795 68.925 282.055 69.015 ;
        RECT 282.315 68.925 282.455 72.580 ;
        RECT 282.775 69.550 282.915 86.125 ;
        RECT 283.635 86.035 283.895 86.125 ;
        RECT 283.635 85.355 283.895 85.675 ;
        RECT 283.695 83.635 283.835 85.355 ;
        RECT 283.635 83.315 283.895 83.635 ;
        RECT 283.635 81.275 283.895 81.595 ;
        RECT 283.175 80.595 283.435 80.915 ;
        RECT 283.235 75.475 283.375 80.595 ;
        RECT 283.695 80.235 283.835 81.275 ;
        RECT 283.635 79.915 283.895 80.235 ;
        RECT 283.175 75.155 283.435 75.475 ;
        RECT 283.235 70.035 283.375 75.155 ;
        RECT 283.695 73.435 283.835 79.915 ;
        RECT 284.095 78.215 284.355 78.535 ;
        RECT 284.155 74.795 284.295 78.215 ;
        RECT 284.095 74.475 284.355 74.795 ;
        RECT 284.615 74.195 284.755 96.575 ;
        RECT 285.535 94.855 285.675 99.635 ;
        RECT 285.935 99.295 286.195 99.615 ;
        RECT 285.995 97.575 286.135 99.295 ;
        RECT 285.935 97.255 286.195 97.575 ;
        RECT 285.475 94.535 285.735 94.855 ;
        RECT 286.455 83.150 286.595 99.635 ;
        RECT 286.915 97.575 287.055 102.615 ;
        RECT 287.775 101.335 288.035 101.655 ;
        RECT 287.835 99.955 287.975 101.335 ;
        RECT 287.775 99.635 288.035 99.955 ;
        RECT 287.835 99.275 287.975 99.635 ;
        RECT 287.775 98.955 288.035 99.275 ;
        RECT 286.855 97.255 287.115 97.575 ;
        RECT 287.835 94.175 287.975 98.955 ;
        RECT 288.295 97.915 288.435 109.225 ;
        RECT 288.695 105.415 288.955 105.735 ;
        RECT 288.755 103.015 288.895 105.415 ;
        RECT 290.075 105.075 290.335 105.395 ;
        RECT 288.695 102.695 288.955 103.015 ;
        RECT 288.755 101.995 288.895 102.695 ;
        RECT 288.695 101.675 288.955 101.995 ;
        RECT 288.235 97.595 288.495 97.915 ;
        RECT 288.755 97.315 288.895 101.675 ;
        RECT 288.295 97.175 288.895 97.315 ;
        RECT 287.775 93.855 288.035 94.175 ;
        RECT 288.295 91.455 288.435 97.175 ;
        RECT 288.695 96.575 288.955 96.895 ;
        RECT 288.235 91.135 288.495 91.455 ;
        RECT 286.855 88.755 287.115 89.075 ;
        RECT 286.915 87.035 287.055 88.755 ;
        RECT 287.765 88.220 288.045 88.590 ;
        RECT 286.855 86.715 287.115 87.035 ;
        RECT 287.835 86.015 287.975 88.220 ;
        RECT 287.315 85.695 287.575 86.015 ;
        RECT 287.775 85.695 288.035 86.015 ;
        RECT 286.385 82.780 286.665 83.150 ;
        RECT 286.455 81.595 286.595 82.780 ;
        RECT 286.395 81.275 286.655 81.595 ;
        RECT 285.015 79.575 285.275 79.895 ;
        RECT 285.075 77.855 285.215 79.575 ;
        RECT 287.375 78.535 287.515 85.695 ;
        RECT 287.315 78.215 287.575 78.535 ;
        RECT 285.015 77.535 285.275 77.855 ;
        RECT 288.755 77.175 288.895 96.575 ;
        RECT 289.155 79.575 289.415 79.895 ;
        RECT 288.695 76.855 288.955 77.175 ;
        RECT 286.395 74.475 286.655 74.795 ;
        RECT 287.765 74.620 288.045 74.990 ;
        RECT 288.235 74.815 288.495 75.135 ;
        RECT 284.155 74.055 284.755 74.195 ;
        RECT 285.475 74.135 285.735 74.455 ;
        RECT 283.635 73.115 283.895 73.435 ;
        RECT 283.175 69.715 283.435 70.035 ;
        RECT 282.705 69.180 282.985 69.550 ;
        RECT 281.795 68.785 282.455 68.925 ;
        RECT 281.795 68.695 282.055 68.785 ;
        RECT 282.315 67.995 282.455 68.785 ;
        RECT 282.255 67.675 282.515 67.995 ;
        RECT 282.255 63.595 282.515 63.915 ;
        RECT 281.335 63.255 281.595 63.575 ;
        RECT 280.875 62.235 281.135 62.555 ;
        RECT 278.115 61.895 278.375 62.215 ;
        RECT 281.395 61.955 281.535 63.255 ;
        RECT 282.315 62.555 282.455 63.595 ;
        RECT 282.255 62.235 282.515 62.555 ;
        RECT 276.275 61.555 276.535 61.875 ;
        RECT 280.935 61.815 281.535 61.955 ;
        RECT 279.955 61.215 280.215 61.535 ;
        RECT 280.015 59.155 280.155 61.215 ;
        RECT 280.935 61.195 281.075 61.815 ;
        RECT 282.775 61.535 282.915 69.180 ;
        RECT 283.235 66.975 283.375 69.715 ;
        RECT 283.175 66.655 283.435 66.975 ;
        RECT 282.715 61.215 282.975 61.535 ;
        RECT 280.875 60.875 281.135 61.195 ;
        RECT 281.795 60.875 282.055 61.195 ;
        RECT 280.935 59.155 281.075 60.875 ;
        RECT 281.855 59.155 281.995 60.875 ;
        RECT 279.955 58.835 280.215 59.155 ;
        RECT 280.875 58.835 281.135 59.155 ;
        RECT 281.795 58.835 282.055 59.155 ;
        RECT 262.935 58.495 263.195 58.815 ;
        RECT 263.395 58.495 263.655 58.815 ;
        RECT 274.435 58.495 274.695 58.815 ;
        RECT 276.275 58.495 276.535 58.815 ;
        RECT 282.715 58.555 282.975 58.815 ;
        RECT 284.155 58.555 284.295 74.055 ;
        RECT 285.535 72.755 285.675 74.135 ;
        RECT 285.475 72.435 285.735 72.755 ;
        RECT 286.455 70.715 286.595 74.475 ;
        RECT 286.855 72.435 287.115 72.755 ;
        RECT 285.935 70.395 286.195 70.715 ;
        RECT 286.395 70.395 286.655 70.715 ;
        RECT 284.555 67.675 284.815 67.995 ;
        RECT 284.615 61.535 284.755 67.675 ;
        RECT 285.995 67.655 286.135 70.395 ;
        RECT 286.915 69.355 287.055 72.435 ;
        RECT 287.835 70.035 287.975 74.620 ;
        RECT 287.775 69.715 288.035 70.035 ;
        RECT 286.855 69.035 287.115 69.355 ;
        RECT 285.935 67.335 286.195 67.655 ;
        RECT 287.775 66.150 288.035 66.295 ;
        RECT 287.765 65.780 288.045 66.150 ;
        RECT 286.855 63.595 287.115 63.915 ;
        RECT 284.555 61.390 284.815 61.535 ;
        RECT 284.545 61.020 284.825 61.390 ;
        RECT 284.555 60.535 284.815 60.855 ;
        RECT 282.715 58.495 284.295 58.555 ;
        RECT 262.995 56.775 263.135 58.495 ;
        RECT 264.315 57.815 264.575 58.135 ;
        RECT 262.935 56.455 263.195 56.775 ;
        RECT 262.475 55.435 262.735 55.755 ;
        RECT 263.395 55.435 263.655 55.755 ;
        RECT 263.455 55.155 263.595 55.435 ;
        RECT 261.155 55.015 263.595 55.155 ;
        RECT 262.935 54.075 263.195 54.395 ;
        RECT 262.995 53.035 263.135 54.075 ;
        RECT 264.375 54.055 264.515 57.815 ;
        RECT 267.995 56.795 268.255 57.115 ;
        RECT 264.775 56.115 265.035 56.435 ;
        RECT 264.315 53.735 264.575 54.055 ;
        RECT 264.835 53.285 264.975 56.115 ;
        RECT 268.055 53.375 268.195 56.795 ;
        RECT 276.335 56.775 276.475 58.495 ;
        RECT 280.875 58.155 281.135 58.475 ;
        RECT 282.775 58.415 284.295 58.495 ;
        RECT 284.615 58.475 284.755 60.535 ;
        RECT 286.915 58.475 287.055 63.595 ;
        RECT 287.835 61.875 287.975 65.780 ;
        RECT 287.775 61.555 288.035 61.875 ;
        RECT 287.835 59.835 287.975 61.555 ;
        RECT 287.775 59.515 288.035 59.835 ;
        RECT 276.735 57.815 276.995 58.135 ;
        RECT 280.935 57.875 281.075 58.155 ;
        RECT 276.795 56.775 276.935 57.815 ;
        RECT 279.095 57.735 281.075 57.875 ;
        RECT 283.635 57.815 283.895 58.135 ;
        RECT 278.575 56.795 278.835 57.115 ;
        RECT 276.275 56.455 276.535 56.775 ;
        RECT 276.735 56.455 276.995 56.775 ;
        RECT 278.115 56.455 278.375 56.775 ;
        RECT 275.355 55.775 275.615 56.095 ;
        RECT 269.375 55.095 269.635 55.415 ;
        RECT 269.435 53.375 269.575 55.095 ;
        RECT 275.415 53.715 275.555 55.775 ;
        RECT 275.355 53.395 275.615 53.715 ;
        RECT 264.375 53.145 264.975 53.285 ;
        RECT 262.935 52.715 263.195 53.035 ;
        RECT 260.635 51.355 260.895 51.675 ;
        RECT 259.245 50.140 259.525 50.510 ;
        RECT 259.315 45.555 259.455 50.140 ;
        RECT 260.175 49.655 260.435 49.975 ;
        RECT 260.235 48.275 260.375 49.655 ;
        RECT 264.375 48.275 264.515 53.145 ;
        RECT 266.615 53.055 266.875 53.375 ;
        RECT 267.535 53.055 267.795 53.375 ;
        RECT 267.995 53.055 268.255 53.375 ;
        RECT 269.375 53.055 269.635 53.375 ;
        RECT 266.675 51.675 266.815 53.055 ;
        RECT 266.615 51.355 266.875 51.675 ;
        RECT 267.595 48.955 267.735 53.055 ;
        RECT 266.615 48.635 266.875 48.955 ;
        RECT 267.535 48.635 267.795 48.955 ;
        RECT 260.175 47.955 260.435 48.275 ;
        RECT 264.315 47.955 264.575 48.275 ;
        RECT 260.235 45.555 260.375 47.955 ;
        RECT 259.255 45.235 259.515 45.555 ;
        RECT 260.175 45.235 260.435 45.555 ;
        RECT 258.795 42.175 259.055 42.495 ;
        RECT 259.255 42.175 259.515 42.495 ;
        RECT 262.935 42.175 263.195 42.495 ;
        RECT 256.955 41.835 257.215 42.155 ;
        RECT 258.335 41.495 258.595 41.815 ;
        RECT 258.395 40.115 258.535 41.495 ;
        RECT 258.335 39.795 258.595 40.115 ;
        RECT 258.795 39.795 259.055 40.115 ;
        RECT 258.395 39.435 258.535 39.795 ;
        RECT 258.335 39.115 258.595 39.435 ;
        RECT 256.955 38.775 257.215 39.095 ;
        RECT 257.415 38.775 257.675 39.095 ;
        RECT 256.035 37.075 256.295 37.395 ;
        RECT 255.115 36.055 255.375 36.375 ;
        RECT 255.175 35.355 255.315 36.055 ;
        RECT 252.355 35.035 252.615 35.355 ;
        RECT 255.115 35.035 255.375 35.355 ;
        RECT 256.095 35.015 256.235 37.075 ;
        RECT 257.015 36.715 257.155 38.775 ;
        RECT 256.955 36.395 257.215 36.715 ;
        RECT 245.055 34.615 246.115 34.755 ;
        RECT 256.035 34.695 256.295 35.015 ;
        RECT 245.055 34.335 245.195 34.615 ;
        RECT 248.215 34.355 248.475 34.675 ;
        RECT 244.995 34.015 245.255 34.335 ;
        RECT 244.535 33.335 244.795 33.655 ;
        RECT 244.595 31.955 244.735 33.335 ;
        RECT 248.275 31.955 248.415 34.355 ;
        RECT 257.475 34.335 257.615 38.775 ;
        RECT 257.415 34.015 257.675 34.335 ;
        RECT 244.535 31.635 244.795 31.955 ;
        RECT 248.215 31.635 248.475 31.955 ;
        RECT 258.855 31.615 258.995 39.795 ;
        RECT 259.315 36.375 259.455 42.175 ;
        RECT 262.475 40.135 262.735 40.455 ;
        RECT 262.015 39.795 262.275 40.115 ;
        RECT 259.255 36.055 259.515 36.375 ;
        RECT 258.795 31.295 259.055 31.615 ;
        RECT 259.315 31.525 259.455 36.055 ;
        RECT 262.075 31.955 262.215 39.795 ;
        RECT 262.535 37.735 262.675 40.135 ;
        RECT 262.995 38.075 263.135 42.175 ;
        RECT 264.375 42.155 264.515 47.955 ;
        RECT 265.235 47.275 265.495 47.595 ;
        RECT 265.295 45.895 265.435 47.275 ;
        RECT 266.675 45.895 266.815 48.635 ;
        RECT 267.535 47.955 267.795 48.275 ;
        RECT 267.595 45.895 267.735 47.955 ;
        RECT 268.915 47.505 269.175 47.595 ;
        RECT 269.435 47.505 269.575 53.055 ;
        RECT 270.755 52.375 271.015 52.695 ;
        RECT 270.815 51.335 270.955 52.375 ;
        RECT 270.755 51.015 271.015 51.335 ;
        RECT 275.415 49.975 275.555 53.395 ;
        RECT 278.175 53.035 278.315 56.455 ;
        RECT 278.635 53.910 278.775 56.795 ;
        RECT 279.095 56.775 279.235 57.735 ;
        RECT 279.035 56.455 279.295 56.775 ;
        RECT 283.695 56.435 283.835 57.815 ;
        RECT 284.155 57.115 284.295 58.415 ;
        RECT 284.555 58.155 284.815 58.475 ;
        RECT 286.855 58.155 287.115 58.475 ;
        RECT 284.095 56.795 284.355 57.115 ;
        RECT 283.635 56.115 283.895 56.435 ;
        RECT 284.155 56.095 284.295 56.795 ;
        RECT 288.295 56.775 288.435 74.815 ;
        RECT 288.755 65.275 288.895 76.855 ;
        RECT 289.215 74.195 289.355 79.575 ;
        RECT 289.615 78.215 289.875 78.535 ;
        RECT 289.675 75.135 289.815 78.215 ;
        RECT 289.615 74.815 289.875 75.135 ;
        RECT 289.615 74.195 289.875 74.455 ;
        RECT 289.215 74.135 289.875 74.195 ;
        RECT 289.215 74.055 289.815 74.135 ;
        RECT 289.675 67.995 289.815 74.055 ;
        RECT 290.135 70.230 290.275 105.075 ;
        RECT 290.595 92.475 290.735 109.225 ;
        RECT 292.375 105.075 292.635 105.395 ;
        RECT 290.535 92.155 290.795 92.475 ;
        RECT 292.435 81.255 292.575 105.075 ;
        RECT 292.895 98.935 293.035 109.225 ;
        RECT 295.195 108.875 295.335 109.225 ;
        RECT 295.655 108.875 295.795 109.415 ;
        RECT 295.195 108.735 295.795 108.875 ;
        RECT 294.675 104.795 294.935 105.055 ;
        RECT 294.675 104.735 295.335 104.795 ;
        RECT 294.735 104.655 295.335 104.735 ;
        RECT 295.195 102.675 295.335 104.655 ;
        RECT 294.675 102.355 294.935 102.675 ;
        RECT 295.135 102.355 295.395 102.675 ;
        RECT 293.755 101.675 294.015 101.995 ;
        RECT 293.815 100.635 293.955 101.675 ;
        RECT 293.755 100.315 294.015 100.635 ;
        RECT 294.735 99.955 294.875 102.355 ;
        RECT 294.675 99.635 294.935 99.955 ;
        RECT 293.755 99.295 294.015 99.615 ;
        RECT 294.215 99.295 294.475 99.615 ;
        RECT 292.835 98.615 293.095 98.935 ;
        RECT 292.835 96.575 293.095 96.895 ;
        RECT 293.815 96.750 293.955 99.295 ;
        RECT 294.275 97.915 294.415 99.295 ;
        RECT 294.215 97.595 294.475 97.915 ;
        RECT 294.275 97.235 294.415 97.595 ;
        RECT 294.735 97.235 294.875 99.635 ;
        RECT 294.215 96.915 294.475 97.235 ;
        RECT 294.675 96.915 294.935 97.235 ;
        RECT 292.375 80.935 292.635 81.255 ;
        RECT 290.995 80.595 291.255 80.915 ;
        RECT 290.535 77.875 290.795 78.195 ;
        RECT 290.595 75.475 290.735 77.875 ;
        RECT 290.535 75.155 290.795 75.475 ;
        RECT 290.595 73.095 290.735 75.155 ;
        RECT 290.535 72.775 290.795 73.095 ;
        RECT 291.055 72.270 291.195 80.595 ;
        RECT 291.915 80.255 292.175 80.575 ;
        RECT 290.985 71.900 291.265 72.270 ;
        RECT 291.055 71.735 291.195 71.900 ;
        RECT 290.995 71.415 291.255 71.735 ;
        RECT 290.065 69.860 290.345 70.230 ;
        RECT 291.975 69.015 292.115 80.255 ;
        RECT 292.375 79.575 292.635 79.895 ;
        RECT 292.435 78.875 292.575 79.575 ;
        RECT 292.375 78.555 292.635 78.875 ;
        RECT 292.435 76.155 292.575 78.555 ;
        RECT 292.375 75.835 292.635 76.155 ;
        RECT 290.075 68.695 290.335 69.015 ;
        RECT 291.915 68.695 292.175 69.015 ;
        RECT 289.615 67.675 289.875 67.995 ;
        RECT 289.675 66.975 289.815 67.675 ;
        RECT 289.615 66.655 289.875 66.975 ;
        RECT 288.695 64.955 288.955 65.275 ;
        RECT 288.755 62.555 288.895 64.955 ;
        RECT 290.135 63.575 290.275 68.695 ;
        RECT 291.975 67.315 292.115 68.695 ;
        RECT 291.915 66.995 292.175 67.315 ;
        RECT 290.075 63.255 290.335 63.575 ;
        RECT 288.695 62.235 288.955 62.555 ;
        RECT 289.615 61.215 289.875 61.535 ;
        RECT 289.675 56.775 289.815 61.215 ;
        RECT 290.535 58.835 290.795 59.155 ;
        RECT 288.235 56.455 288.495 56.775 ;
        RECT 289.615 56.455 289.875 56.775 ;
        RECT 284.095 55.775 284.355 56.095 ;
        RECT 285.935 55.775 286.195 56.095 ;
        RECT 278.565 53.540 278.845 53.910 ;
        RECT 280.415 53.735 280.675 54.055 ;
        RECT 278.115 52.715 278.375 53.035 ;
        RECT 276.735 51.355 276.995 51.675 ;
        RECT 271.675 49.655 271.935 49.975 ;
        RECT 275.355 49.655 275.615 49.975 ;
        RECT 268.915 47.365 269.575 47.505 ;
        RECT 268.915 47.275 269.175 47.365 ;
        RECT 265.235 45.575 265.495 45.895 ;
        RECT 266.615 45.575 266.875 45.895 ;
        RECT 267.535 45.575 267.795 45.895 ;
        RECT 264.775 44.555 265.035 44.875 ;
        RECT 264.315 41.835 264.575 42.155 ;
        RECT 264.835 40.795 264.975 44.555 ;
        RECT 265.295 42.155 265.435 45.575 ;
        RECT 268.975 45.555 269.115 47.275 ;
        RECT 268.915 45.235 269.175 45.555 ;
        RECT 267.535 44.215 267.795 44.535 ;
        RECT 267.595 42.835 267.735 44.215 ;
        RECT 267.535 42.515 267.795 42.835 ;
        RECT 265.235 41.835 265.495 42.155 ;
        RECT 264.775 40.475 265.035 40.795 ;
        RECT 268.975 40.455 269.115 45.235 ;
        RECT 269.835 44.895 270.095 45.215 ;
        RECT 269.895 43.515 270.035 44.895 ;
        RECT 270.755 44.215 271.015 44.535 ;
        RECT 269.835 43.195 270.095 43.515 ;
        RECT 270.815 41.815 270.955 44.215 ;
        RECT 270.755 41.495 271.015 41.815 ;
        RECT 268.915 40.135 269.175 40.455 ;
        RECT 267.075 39.455 267.335 39.775 ;
        RECT 266.615 38.775 266.875 39.095 ;
        RECT 262.935 37.755 263.195 38.075 ;
        RECT 262.475 37.415 262.735 37.735 ;
        RECT 262.995 37.055 263.135 37.755 ;
        RECT 266.675 37.055 266.815 38.775 ;
        RECT 267.135 37.055 267.275 39.455 ;
        RECT 268.975 39.095 269.115 40.135 ;
        RECT 270.815 39.095 270.955 41.495 ;
        RECT 268.915 38.775 269.175 39.095 ;
        RECT 270.755 38.775 271.015 39.095 ;
        RECT 262.935 36.735 263.195 37.055 ;
        RECT 266.615 36.735 266.875 37.055 ;
        RECT 267.075 36.735 267.335 37.055 ;
        RECT 267.135 35.355 267.275 36.735 ;
        RECT 267.075 35.035 267.335 35.355 ;
        RECT 271.735 34.675 271.875 49.655 ;
        RECT 273.055 47.615 273.315 47.935 ;
        RECT 273.115 46.235 273.255 47.615 ;
        RECT 273.055 45.915 273.315 46.235 ;
        RECT 272.135 45.235 272.395 45.555 ;
        RECT 272.195 40.705 272.335 45.235 ;
        RECT 274.435 44.895 274.695 45.215 ;
        RECT 274.495 43.515 274.635 44.895 ;
        RECT 274.435 43.195 274.695 43.515 ;
        RECT 276.795 42.155 276.935 51.355 ;
        RECT 278.175 51.335 278.315 52.715 ;
        RECT 278.635 52.695 278.775 53.540 ;
        RECT 278.575 52.375 278.835 52.695 ;
        RECT 278.115 51.015 278.375 51.335 ;
        RECT 279.035 49.995 279.295 50.315 ;
        RECT 279.095 45.555 279.235 49.995 ;
        RECT 279.495 49.655 279.755 49.975 ;
        RECT 279.555 48.275 279.695 49.655 ;
        RECT 279.495 47.955 279.755 48.275 ;
        RECT 280.475 47.935 280.615 53.735 ;
        RECT 285.995 53.715 286.135 55.775 ;
        RECT 288.295 54.395 288.435 56.455 ;
        RECT 288.235 54.075 288.495 54.395 ;
        RECT 285.935 53.395 286.195 53.715 ;
        RECT 285.995 50.655 286.135 53.395 ;
        RECT 288.295 53.375 288.435 54.075 ;
        RECT 290.595 53.715 290.735 58.835 ;
        RECT 292.895 57.115 293.035 96.575 ;
        RECT 293.745 96.380 294.025 96.750 ;
        RECT 293.815 95.195 293.955 96.380 ;
        RECT 293.755 94.875 294.015 95.195 ;
        RECT 293.295 94.195 293.555 94.515 ;
        RECT 293.355 91.795 293.495 94.195 ;
        RECT 293.755 93.175 294.015 93.495 ;
        RECT 293.815 91.795 293.955 93.175 ;
        RECT 293.295 91.475 293.555 91.795 ;
        RECT 293.755 91.475 294.015 91.795 ;
        RECT 293.355 89.755 293.495 91.475 ;
        RECT 295.195 91.455 295.335 102.355 ;
        RECT 296.515 101.335 296.775 101.655 ;
        RECT 296.055 96.915 296.315 97.235 ;
        RECT 295.595 94.535 295.855 94.855 ;
        RECT 295.135 91.365 295.395 91.455 ;
        RECT 294.735 91.225 295.395 91.365 ;
        RECT 293.295 89.435 293.555 89.755 ;
        RECT 294.735 88.735 294.875 91.225 ;
        RECT 295.135 91.135 295.395 91.225 ;
        RECT 294.675 88.415 294.935 88.735 ;
        RECT 294.735 86.015 294.875 88.415 ;
        RECT 294.675 85.695 294.935 86.015 ;
        RECT 295.655 85.675 295.795 94.535 ;
        RECT 295.595 85.355 295.855 85.675 ;
        RECT 296.115 83.635 296.255 96.915 ;
        RECT 296.575 96.555 296.715 101.335 ;
        RECT 296.515 96.235 296.775 96.555 ;
        RECT 297.035 95.955 297.175 109.415 ;
        RECT 297.425 109.225 297.705 141.105 ;
        RECT 299.725 109.225 300.005 141.685 ;
        RECT 302.025 109.225 302.305 142.265 ;
        RECT 304.325 109.225 304.605 142.845 ;
        RECT 306.625 109.225 306.905 143.425 ;
        RECT 308.925 109.225 309.205 144.005 ;
        RECT 296.575 95.815 297.175 95.955 ;
        RECT 296.575 92.135 296.715 95.815 ;
        RECT 296.975 94.875 297.235 95.195 ;
        RECT 296.515 91.815 296.775 92.135 ;
        RECT 296.515 90.455 296.775 90.775 ;
        RECT 296.575 89.415 296.715 90.455 ;
        RECT 296.515 89.095 296.775 89.415 ;
        RECT 297.035 83.975 297.175 94.875 ;
        RECT 297.495 87.115 297.635 109.225 ;
        RECT 298.355 105.645 298.615 105.735 ;
        RECT 298.355 105.505 299.015 105.645 ;
        RECT 298.355 105.415 298.615 105.505 ;
        RECT 297.895 102.355 298.155 102.675 ;
        RECT 297.955 97.915 298.095 102.355 ;
        RECT 298.355 101.335 298.615 101.655 ;
        RECT 298.415 100.635 298.555 101.335 ;
        RECT 298.355 100.315 298.615 100.635 ;
        RECT 298.415 97.915 298.555 100.315 ;
        RECT 298.875 100.295 299.015 105.505 ;
        RECT 299.275 101.335 299.535 101.655 ;
        RECT 299.335 100.830 299.475 101.335 ;
        RECT 299.265 100.460 299.545 100.830 ;
        RECT 299.795 100.545 299.935 109.225 ;
        RECT 302.095 106.155 302.235 109.225 ;
        RECT 302.095 106.075 302.695 106.155 ;
        RECT 302.095 106.015 302.755 106.075 ;
        RECT 302.495 105.755 302.755 106.015 ;
        RECT 303.415 105.075 303.675 105.395 ;
        RECT 303.475 104.375 303.615 105.075 ;
        RECT 303.875 104.735 304.135 105.055 ;
        RECT 303.415 104.055 303.675 104.375 ;
        RECT 303.475 102.335 303.615 104.055 ;
        RECT 303.935 103.355 304.075 104.735 ;
        RECT 303.875 103.035 304.135 103.355 ;
        RECT 302.495 102.015 302.755 102.335 ;
        RECT 303.415 102.015 303.675 102.335 ;
        RECT 300.655 100.545 300.915 100.635 ;
        RECT 298.815 99.975 299.075 100.295 ;
        RECT 297.895 97.595 298.155 97.915 ;
        RECT 298.355 97.595 298.615 97.915 ;
        RECT 297.955 95.275 298.095 97.595 ;
        RECT 298.875 96.070 299.015 99.975 ;
        RECT 298.805 95.700 299.085 96.070 ;
        RECT 297.955 95.135 298.555 95.275 ;
        RECT 297.885 94.340 298.165 94.710 ;
        RECT 297.955 91.455 298.095 94.340 ;
        RECT 298.415 93.495 298.555 95.135 ;
        RECT 298.805 95.020 299.085 95.390 ;
        RECT 298.815 94.875 299.075 95.020 ;
        RECT 298.355 93.175 298.615 93.495 ;
        RECT 299.335 91.875 299.475 100.460 ;
        RECT 299.795 100.405 300.915 100.545 ;
        RECT 300.655 100.315 300.915 100.405 ;
        RECT 301.115 99.295 301.375 99.615 ;
        RECT 301.175 97.575 301.315 99.295 ;
        RECT 301.115 97.255 301.375 97.575 ;
        RECT 299.735 96.915 299.995 97.235 ;
        RECT 299.795 94.175 299.935 96.915 ;
        RECT 300.185 95.700 300.465 96.070 ;
        RECT 299.735 93.855 299.995 94.175 ;
        RECT 298.875 91.795 299.475 91.875 ;
        RECT 299.795 91.795 299.935 93.855 ;
        RECT 298.815 91.735 299.475 91.795 ;
        RECT 298.815 91.475 299.075 91.735 ;
        RECT 299.735 91.475 299.995 91.795 ;
        RECT 297.895 91.365 298.155 91.455 ;
        RECT 297.895 91.225 298.555 91.365 ;
        RECT 297.895 91.135 298.155 91.225 ;
        RECT 298.415 88.735 298.555 91.225 ;
        RECT 298.815 90.795 299.075 91.115 ;
        RECT 298.355 88.415 298.615 88.735 ;
        RECT 297.495 87.035 298.095 87.115 ;
        RECT 297.495 86.975 298.155 87.035 ;
        RECT 297.895 86.715 298.155 86.975 ;
        RECT 296.975 83.655 297.235 83.975 ;
        RECT 295.135 83.315 295.395 83.635 ;
        RECT 296.055 83.315 296.315 83.635 ;
        RECT 294.675 80.935 294.935 81.255 ;
        RECT 294.215 79.575 294.475 79.895 ;
        RECT 294.275 74.795 294.415 79.575 ;
        RECT 294.735 77.175 294.875 80.935 ;
        RECT 295.195 77.855 295.335 83.315 ;
        RECT 296.115 80.915 296.255 83.315 ;
        RECT 296.055 80.595 296.315 80.915 ;
        RECT 296.115 78.195 296.255 80.595 ;
        RECT 296.055 77.875 296.315 78.195 ;
        RECT 295.135 77.535 295.395 77.855 ;
        RECT 294.675 76.855 294.935 77.175 ;
        RECT 294.675 75.045 294.935 75.135 ;
        RECT 295.195 75.045 295.335 77.535 ;
        RECT 298.355 75.155 298.615 75.475 ;
        RECT 294.675 74.905 295.335 75.045 ;
        RECT 294.675 74.815 294.935 74.905 ;
        RECT 294.215 74.475 294.475 74.795 ;
        RECT 293.285 72.580 293.565 72.950 ;
        RECT 293.355 71.735 293.495 72.580 ;
        RECT 294.735 72.415 294.875 74.815 ;
        RECT 298.415 73.095 298.555 75.155 ;
        RECT 298.355 72.775 298.615 73.095 ;
        RECT 294.675 72.095 294.935 72.415 ;
        RECT 293.295 71.415 293.555 71.735 ;
        RECT 293.355 70.230 293.495 71.415 ;
        RECT 293.285 69.860 293.565 70.230 ;
        RECT 294.215 69.605 294.475 69.695 ;
        RECT 294.735 69.605 294.875 72.095 ;
        RECT 295.595 71.415 295.855 71.735 ;
        RECT 294.215 69.465 294.875 69.605 ;
        RECT 294.215 69.375 294.475 69.465 ;
        RECT 294.275 65.275 294.415 69.375 ;
        RECT 295.655 66.715 295.795 71.415 ;
        RECT 296.055 69.035 296.315 69.355 ;
        RECT 296.115 67.995 296.255 69.035 ;
        RECT 296.055 67.675 296.315 67.995 ;
        RECT 298.355 66.995 298.615 67.315 ;
        RECT 296.045 66.715 296.325 66.830 ;
        RECT 295.655 66.575 296.325 66.715 ;
        RECT 296.045 66.460 296.325 66.575 ;
        RECT 294.215 64.955 294.475 65.275 ;
        RECT 294.275 64.595 294.415 64.955 ;
        RECT 294.215 64.275 294.475 64.595 ;
        RECT 295.135 63.595 295.395 63.915 ;
        RECT 295.195 62.555 295.335 63.595 ;
        RECT 296.115 62.555 296.255 66.460 ;
        RECT 296.975 66.315 297.235 66.635 ;
        RECT 297.035 64.675 297.175 66.315 ;
        RECT 297.035 64.595 297.635 64.675 ;
        RECT 297.035 64.535 297.695 64.595 ;
        RECT 296.515 63.255 296.775 63.575 ;
        RECT 295.135 62.235 295.395 62.555 ;
        RECT 296.055 62.235 296.315 62.555 ;
        RECT 293.755 59.175 294.015 59.495 ;
        RECT 293.815 58.135 293.955 59.175 ;
        RECT 293.755 57.815 294.015 58.135 ;
        RECT 292.835 56.795 293.095 57.115 ;
        RECT 293.815 56.435 293.955 57.815 ;
        RECT 296.115 57.115 296.255 62.235 ;
        RECT 296.575 62.215 296.715 63.255 ;
        RECT 296.515 62.070 296.775 62.215 ;
        RECT 296.505 61.700 296.785 62.070 ;
        RECT 297.035 61.195 297.175 64.535 ;
        RECT 297.435 64.275 297.695 64.535 ;
        RECT 297.895 63.595 298.155 63.915 ;
        RECT 296.975 60.875 297.235 61.195 ;
        RECT 297.955 58.135 298.095 63.595 ;
        RECT 298.415 61.535 298.555 66.995 ;
        RECT 298.875 66.295 299.015 90.795 ;
        RECT 300.255 90.775 300.395 95.700 ;
        RECT 302.025 95.020 302.305 95.390 ;
        RECT 300.195 90.455 300.455 90.775 ;
        RECT 300.255 89.415 300.395 90.455 ;
        RECT 300.195 89.095 300.455 89.415 ;
        RECT 299.735 85.585 299.995 85.675 ;
        RECT 300.255 85.585 300.395 89.095 ;
        RECT 302.095 88.055 302.235 95.020 ;
        RECT 302.555 94.515 302.695 102.015 ;
        RECT 302.955 98.955 303.215 99.275 ;
        RECT 303.015 95.390 303.155 98.955 ;
        RECT 303.475 97.430 303.615 102.015 ;
        RECT 303.875 99.975 304.135 100.295 ;
        RECT 304.395 100.035 304.535 109.225 ;
        RECT 304.795 106.775 305.055 107.095 ;
        RECT 304.855 104.715 304.995 106.775 ;
        RECT 304.795 104.395 305.055 104.715 ;
        RECT 305.255 102.695 305.515 103.015 ;
        RECT 303.405 97.060 303.685 97.430 ;
        RECT 302.945 95.020 303.225 95.390 ;
        RECT 303.415 94.535 303.675 94.855 ;
        RECT 302.495 94.195 302.755 94.515 ;
        RECT 302.555 91.875 302.695 94.195 ;
        RECT 302.555 91.735 303.155 91.875 ;
        RECT 302.495 90.795 302.755 91.115 ;
        RECT 302.035 87.735 302.295 88.055 ;
        RECT 299.735 85.445 300.395 85.585 ;
        RECT 299.735 85.355 299.995 85.445 ;
        RECT 299.795 83.975 299.935 85.355 ;
        RECT 302.095 84.315 302.235 87.735 ;
        RECT 302.035 83.995 302.295 84.315 ;
        RECT 299.735 83.655 299.995 83.975 ;
        RECT 302.555 79.895 302.695 90.795 ;
        RECT 303.015 85.335 303.155 91.735 ;
        RECT 302.955 85.015 303.215 85.335 ;
        RECT 302.495 79.575 302.755 79.895 ;
        RECT 302.555 78.535 302.695 79.575 ;
        RECT 302.495 78.215 302.755 78.535 ;
        RECT 302.555 74.795 302.695 78.215 ;
        RECT 302.955 76.855 303.215 77.175 ;
        RECT 303.015 75.135 303.155 76.855 ;
        RECT 302.955 74.815 303.215 75.135 ;
        RECT 302.495 74.475 302.755 74.795 ;
        RECT 302.955 73.115 303.215 73.435 ;
        RECT 303.475 73.395 303.615 94.535 ;
        RECT 303.935 88.735 304.075 99.975 ;
        RECT 304.395 99.895 304.995 100.035 ;
        RECT 304.855 95.195 304.995 99.895 ;
        RECT 305.315 96.895 305.455 102.695 ;
        RECT 305.715 98.675 305.975 98.935 ;
        RECT 305.715 98.615 306.375 98.675 ;
        RECT 305.775 98.535 306.375 98.615 ;
        RECT 305.255 96.575 305.515 96.895 ;
        RECT 304.795 94.875 305.055 95.195 ;
        RECT 303.875 88.415 304.135 88.735 ;
        RECT 304.335 79.915 304.595 80.235 ;
        RECT 304.395 76.155 304.535 79.915 ;
        RECT 304.795 77.195 305.055 77.515 ;
        RECT 304.335 75.835 304.595 76.155 ;
        RECT 303.475 73.255 304.075 73.395 ;
        RECT 299.275 72.775 299.535 73.095 ;
        RECT 303.015 72.950 303.155 73.115 ;
        RECT 299.335 69.015 299.475 72.775 ;
        RECT 302.945 72.580 303.225 72.950 ;
        RECT 303.415 72.270 303.675 72.415 ;
        RECT 303.405 71.900 303.685 72.270 ;
        RECT 302.495 69.035 302.755 69.355 ;
        RECT 299.275 68.695 299.535 69.015 ;
        RECT 299.275 66.655 299.535 66.975 ;
        RECT 300.655 66.655 300.915 66.975 ;
        RECT 298.815 65.975 299.075 66.295 ;
        RECT 299.335 65.275 299.475 66.655 ;
        RECT 300.715 65.275 300.855 66.655 ;
        RECT 299.275 64.955 299.535 65.275 ;
        RECT 300.655 64.955 300.915 65.275 ;
        RECT 302.555 62.215 302.695 69.035 ;
        RECT 303.935 69.015 304.075 73.255 ;
        RECT 304.855 70.715 304.995 77.195 ;
        RECT 305.315 71.735 305.455 96.575 ;
        RECT 306.235 96.215 306.375 98.535 ;
        RECT 306.175 95.895 306.435 96.215 ;
        RECT 305.715 94.195 305.975 94.515 ;
        RECT 305.255 71.415 305.515 71.735 ;
        RECT 304.795 70.395 305.055 70.715 ;
        RECT 303.875 68.695 304.135 69.015 ;
        RECT 303.935 67.995 304.075 68.695 ;
        RECT 303.875 67.675 304.135 67.995 ;
        RECT 304.335 67.335 304.595 67.655 ;
        RECT 302.495 61.895 302.755 62.215 ;
        RECT 301.115 61.555 301.375 61.875 ;
        RECT 298.355 61.215 298.615 61.535 ;
        RECT 301.175 59.835 301.315 61.555 ;
        RECT 302.035 60.535 302.295 60.855 ;
        RECT 301.115 59.515 301.375 59.835 ;
        RECT 302.095 58.475 302.235 60.535 ;
        RECT 302.035 58.155 302.295 58.475 ;
        RECT 297.895 57.815 298.155 58.135 ;
        RECT 296.055 56.795 296.315 57.115 ;
        RECT 297.955 56.775 298.095 57.815 ;
        RECT 297.895 56.455 298.155 56.775 ;
        RECT 293.755 56.115 294.015 56.435 ;
        RECT 291.455 55.095 291.715 55.415 ;
        RECT 290.535 53.395 290.795 53.715 ;
        RECT 288.235 53.055 288.495 53.375 ;
        RECT 290.595 50.995 290.735 53.395 ;
        RECT 291.515 53.035 291.655 55.095 ;
        RECT 297.955 54.395 298.095 56.455 ;
        RECT 297.895 54.075 298.155 54.395 ;
        RECT 291.915 53.735 292.175 54.055 ;
        RECT 291.455 52.715 291.715 53.035 ;
        RECT 290.535 50.675 290.795 50.995 ;
        RECT 285.935 50.335 286.195 50.655 ;
        RECT 286.855 50.335 287.115 50.655 ;
        RECT 280.415 47.615 280.675 47.935 ;
        RECT 280.475 46.235 280.615 47.615 ;
        RECT 280.415 45.915 280.675 46.235 ;
        RECT 279.035 45.235 279.295 45.555 ;
        RECT 285.995 45.215 286.135 50.335 ;
        RECT 286.915 48.955 287.055 50.335 ;
        RECT 286.855 48.635 287.115 48.955 ;
        RECT 290.595 48.615 290.735 50.675 ;
        RECT 290.535 48.295 290.795 48.615 ;
        RECT 285.475 44.895 285.735 45.215 ;
        RECT 285.935 44.895 286.195 45.215 ;
        RECT 281.335 42.175 281.595 42.495 ;
        RECT 276.735 41.835 276.995 42.155 ;
        RECT 277.655 41.495 277.915 41.815 ;
        RECT 278.115 41.495 278.375 41.815 ;
        RECT 273.055 40.705 273.315 40.795 ;
        RECT 272.195 40.565 273.315 40.705 ;
        RECT 272.195 39.775 272.335 40.565 ;
        RECT 273.055 40.475 273.315 40.565 ;
        RECT 277.715 40.115 277.855 41.495 ;
        RECT 276.275 39.795 276.535 40.115 ;
        RECT 277.655 39.795 277.915 40.115 ;
        RECT 272.135 39.455 272.395 39.775 ;
        RECT 276.335 39.515 276.475 39.795 ;
        RECT 276.335 39.375 276.935 39.515 ;
        RECT 273.055 38.775 273.315 39.095 ;
        RECT 273.115 35.015 273.255 38.775 ;
        RECT 276.795 38.075 276.935 39.375 ;
        RECT 276.735 37.755 276.995 38.075 ;
        RECT 278.175 37.395 278.315 41.495 ;
        RECT 281.395 40.795 281.535 42.175 ;
        RECT 281.335 40.705 281.595 40.795 ;
        RECT 280.935 40.565 281.595 40.705 ;
        RECT 280.415 37.755 280.675 38.075 ;
        RECT 278.115 37.075 278.375 37.395 ;
        RECT 279.495 36.395 279.755 36.715 ;
        RECT 279.555 35.015 279.695 36.395 ;
        RECT 280.475 35.355 280.615 37.755 ;
        RECT 280.935 36.715 281.075 40.565 ;
        RECT 281.335 40.475 281.595 40.565 ;
        RECT 285.535 39.775 285.675 44.895 ;
        RECT 290.595 42.835 290.735 48.295 ;
        RECT 291.455 47.275 291.715 47.595 ;
        RECT 290.535 42.515 290.795 42.835 ;
        RECT 291.515 42.155 291.655 47.275 ;
        RECT 291.975 47.255 292.115 53.735 ;
        RECT 294.215 52.715 294.475 53.035 ;
        RECT 294.275 47.595 294.415 52.715 ;
        RECT 297.955 51.335 298.095 54.075 ;
        RECT 300.195 53.055 300.455 53.375 ;
        RECT 304.395 53.115 304.535 67.335 ;
        RECT 305.315 62.215 305.455 71.415 ;
        RECT 305.775 63.575 305.915 94.195 ;
        RECT 306.235 94.030 306.375 95.895 ;
        RECT 306.695 95.195 306.835 109.225 ;
        RECT 308.475 105.075 308.735 105.395 ;
        RECT 307.095 101.335 307.355 101.655 ;
        RECT 307.155 96.555 307.295 101.335 ;
        RECT 307.095 96.235 307.355 96.555 ;
        RECT 306.635 94.875 306.895 95.195 ;
        RECT 306.165 93.660 306.445 94.030 ;
        RECT 306.235 86.355 306.375 93.660 ;
        RECT 307.095 91.815 307.355 92.135 ;
        RECT 307.155 89.755 307.295 91.815 ;
        RECT 307.095 89.435 307.355 89.755 ;
        RECT 308.015 88.755 308.275 89.075 ;
        RECT 306.175 86.035 306.435 86.355 ;
        RECT 307.555 85.695 307.815 86.015 ;
        RECT 307.615 85.190 307.755 85.695 ;
        RECT 307.545 84.820 307.825 85.190 ;
        RECT 306.635 81.275 306.895 81.595 ;
        RECT 306.695 78.875 306.835 81.275 ;
        RECT 306.635 78.785 306.895 78.875 ;
        RECT 306.235 78.645 306.895 78.785 ;
        RECT 306.235 69.695 306.375 78.645 ;
        RECT 306.635 78.555 306.895 78.645 ;
        RECT 307.095 75.155 307.355 75.475 ;
        RECT 307.155 72.755 307.295 75.155 ;
        RECT 307.095 72.435 307.355 72.755 ;
        RECT 307.555 72.435 307.815 72.755 ;
        RECT 307.155 70.035 307.295 72.435 ;
        RECT 307.095 69.715 307.355 70.035 ;
        RECT 306.175 69.375 306.435 69.695 ;
        RECT 306.635 68.695 306.895 69.015 ;
        RECT 306.695 63.575 306.835 68.695 ;
        RECT 305.715 63.255 305.975 63.575 ;
        RECT 306.635 63.255 306.895 63.575 ;
        RECT 306.695 62.555 306.835 63.255 ;
        RECT 306.635 62.235 306.895 62.555 ;
        RECT 305.255 61.895 305.515 62.215 ;
        RECT 307.615 56.515 307.755 72.435 ;
        RECT 308.075 68.870 308.215 88.755 ;
        RECT 308.535 73.395 308.675 105.075 ;
        RECT 308.995 101.905 309.135 109.225 ;
        RECT 308.995 101.765 309.595 101.905 ;
        RECT 308.925 101.140 309.205 101.510 ;
        RECT 308.995 92.475 309.135 101.140 ;
        RECT 308.935 92.155 309.195 92.475 ;
        RECT 309.455 89.755 309.595 101.765 ;
        RECT 309.855 91.135 310.115 91.455 ;
        RECT 309.395 89.435 309.655 89.755 ;
        RECT 308.535 73.255 309.135 73.395 ;
        RECT 308.005 68.500 308.285 68.870 ;
        RECT 308.475 68.695 308.735 69.015 ;
        RECT 308.075 67.995 308.215 68.500 ;
        RECT 308.015 67.675 308.275 67.995 ;
        RECT 308.075 64.255 308.215 67.675 ;
        RECT 308.015 63.935 308.275 64.255 ;
        RECT 300.255 51.675 300.395 53.055 ;
        RECT 303.935 53.035 304.535 53.115 ;
        RECT 303.875 52.975 304.535 53.035 ;
        RECT 303.875 52.715 304.135 52.975 ;
        RECT 300.195 51.355 300.455 51.675 ;
        RECT 297.895 51.015 298.155 51.335 ;
        RECT 294.215 47.275 294.475 47.595 ;
        RECT 291.915 46.935 292.175 47.255 ;
        RECT 292.835 46.935 293.095 47.255 ;
        RECT 292.895 42.155 293.035 46.935 ;
        RECT 304.395 45.555 304.535 52.975 ;
        RECT 307.155 56.375 307.755 56.515 ;
        RECT 304.335 45.235 304.595 45.555 ;
        RECT 305.255 45.235 305.515 45.555 ;
        RECT 296.515 44.895 296.775 45.215 ;
        RECT 291.455 41.835 291.715 42.155 ;
        RECT 292.835 41.835 293.095 42.155 ;
        RECT 282.715 39.455 282.975 39.775 ;
        RECT 285.475 39.455 285.735 39.775 ;
        RECT 281.335 38.775 281.595 39.095 ;
        RECT 281.395 37.735 281.535 38.775 ;
        RECT 282.775 38.075 282.915 39.455 ;
        RECT 291.515 39.095 291.655 41.835 ;
        RECT 296.575 40.795 296.715 44.895 ;
        RECT 304.395 44.875 304.535 45.235 ;
        RECT 304.335 44.555 304.595 44.875 ;
        RECT 296.515 40.475 296.775 40.795 ;
        RECT 304.395 40.455 304.535 44.555 ;
        RECT 304.795 44.215 305.055 44.535 ;
        RECT 304.855 42.495 304.995 44.215 ;
        RECT 304.795 42.175 305.055 42.495 ;
        RECT 305.315 41.815 305.455 45.235 ;
        RECT 306.175 44.215 306.435 44.535 ;
        RECT 306.235 42.835 306.375 44.215 ;
        RECT 306.175 42.515 306.435 42.835 ;
        RECT 307.155 42.495 307.295 56.375 ;
        RECT 307.555 55.775 307.815 56.095 ;
        RECT 307.615 54.395 307.755 55.775 ;
        RECT 307.555 54.075 307.815 54.395 ;
        RECT 308.535 50.995 308.675 68.695 ;
        RECT 308.995 61.875 309.135 73.255 ;
        RECT 309.395 69.375 309.655 69.695 ;
        RECT 309.455 68.870 309.595 69.375 ;
        RECT 309.385 68.500 309.665 68.870 ;
        RECT 308.935 61.555 309.195 61.875 ;
        RECT 308.935 58.835 309.195 59.155 ;
        RECT 308.995 56.095 309.135 58.835 ;
        RECT 308.935 55.775 309.195 56.095 ;
        RECT 308.995 50.995 309.135 55.775 ;
        RECT 309.395 53.055 309.655 53.375 ;
        RECT 309.455 52.550 309.595 53.055 ;
        RECT 309.385 52.180 309.665 52.550 ;
        RECT 308.475 50.675 308.735 50.995 ;
        RECT 308.935 50.675 309.195 50.995 ;
        RECT 309.915 49.975 310.055 91.135 ;
        RECT 310.315 86.375 310.575 86.695 ;
        RECT 309.855 49.655 310.115 49.975 ;
        RECT 310.375 45.215 310.515 86.375 ;
        RECT 310.315 44.895 310.575 45.215 ;
        RECT 307.095 42.235 307.355 42.495 ;
        RECT 307.095 42.175 307.755 42.235 ;
        RECT 307.155 42.095 307.755 42.175 ;
        RECT 305.255 41.495 305.515 41.815 ;
        RECT 307.095 41.495 307.355 41.815 ;
        RECT 307.155 40.455 307.295 41.495 ;
        RECT 304.335 40.135 304.595 40.455 ;
        RECT 307.095 40.135 307.355 40.455 ;
        RECT 283.175 38.775 283.435 39.095 ;
        RECT 291.455 38.775 291.715 39.095 ;
        RECT 282.715 37.755 282.975 38.075 ;
        RECT 281.335 37.415 281.595 37.735 ;
        RECT 280.875 36.395 281.135 36.715 ;
        RECT 280.415 35.035 280.675 35.355 ;
        RECT 283.235 35.015 283.375 38.775 ;
        RECT 307.615 37.735 307.755 42.095 ;
        RECT 307.555 37.415 307.815 37.735 ;
        RECT 308.935 36.395 309.195 36.715 ;
        RECT 308.995 36.230 309.135 36.395 ;
        RECT 308.925 35.860 309.205 36.230 ;
        RECT 316.555 35.745 318.485 36.545 ;
        RECT 273.055 34.695 273.315 35.015 ;
        RECT 279.495 34.695 279.755 35.015 ;
        RECT 283.175 34.695 283.435 35.015 ;
        RECT 271.675 34.355 271.935 34.675 ;
        RECT 262.015 31.635 262.275 31.955 ;
        RECT 259.715 31.525 259.975 31.615 ;
        RECT 259.315 31.385 259.975 31.525 ;
        RECT 259.715 31.295 259.975 31.385 ;
        RECT 243.615 30.955 243.875 31.275 ;
        RECT 243.155 30.615 243.415 30.935 ;
        RECT 212.335 26.875 212.595 27.195 ;
        RECT 206.815 26.195 207.075 26.515 ;
        RECT 199.915 25.855 200.175 26.175 ;
        RECT 10.170 23.510 74.550 25.010 ;
        RECT 79.810 23.665 127.975 24.765 ;
        RECT 180.945 24.640 182.485 25.010 ;
        RECT 10.170 21.510 74.550 23.010 ;
        RECT 79.810 22.165 127.975 23.265 ;
        RECT 177.645 21.920 179.185 22.290 ;
        RECT 79.810 20.665 127.975 21.765 ;
        RECT 10.170 18.105 74.550 20.485 ;
        RECT 79.810 19.165 127.975 20.265 ;
        RECT 141.295 19.425 143.400 20.015 ;
        RECT 180.945 19.200 182.485 19.570 ;
        RECT 10.170 15.580 74.550 17.080 ;
        RECT 177.645 16.480 179.185 16.850 ;
        RECT 10.170 13.580 74.550 15.080 ;
        RECT 180.945 13.760 182.485 14.130 ;
        RECT 10.170 11.580 74.550 13.080 ;
        RECT 10.170 9.555 74.550 10.555 ;
        RECT 80.745 9.665 82.345 10.465 ;
        RECT 7.065 5.690 8.665 8.890 ;
        RECT 14.965 5.690 16.565 8.890 ;
        RECT 128.965 5.690 130.565 8.890 ;
      LAYER met3 ;
        RECT 125.730 225.710 126.530 225.760 ;
        RECT 23.260 225.160 23.660 225.560 ;
        RECT 1.000 224.760 23.660 225.160 ;
        RECT 45.340 224.760 45.740 225.560 ;
        RECT 64.710 225.310 65.510 225.710 ;
        RECT 125.730 225.410 252.160 225.710 ;
        RECT 125.730 225.360 126.530 225.410 ;
        RECT 59.190 224.760 59.990 225.160 ;
        RECT 1.000 221.560 1.400 224.760 ;
        RECT 67.470 224.710 68.270 225.110 ;
        RECT 129.395 225.050 130.195 225.100 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.110 71.030 224.510 ;
        RECT 72.990 223.510 73.790 223.910 ;
        RECT 75.700 223.310 76.100 224.860 ;
        RECT 75.700 222.910 76.500 223.310 ;
        RECT 78.545 222.710 78.945 224.860 ;
        RECT 78.545 222.310 79.345 222.710 ;
        RECT 83.980 222.110 84.380 224.860 ;
        RECT 83.980 221.710 84.780 222.110 ;
        RECT 1.000 220.760 1.800 221.560 ;
        RECT 86.740 221.510 87.140 224.860 ;
        RECT 86.740 221.110 87.540 221.510 ;
        RECT 92.260 220.910 92.660 224.860 ;
        RECT 129.375 224.750 251.225 225.050 ;
        RECT 129.395 224.700 130.195 224.750 ;
        RECT 108.865 224.515 109.665 224.615 ;
        RECT 95.020 223.650 95.420 224.450 ;
        RECT 97.780 223.650 98.180 224.450 ;
        RECT 100.540 223.650 100.940 224.450 ;
        RECT 103.300 223.650 103.700 224.450 ;
        RECT 106.060 223.915 106.460 224.450 ;
        RECT 108.865 224.215 129.040 224.515 ;
        RECT 95.070 221.515 95.370 223.650 ;
        RECT 97.830 222.115 98.130 223.650 ;
        RECT 100.590 222.715 100.890 223.650 ;
        RECT 103.350 223.315 103.650 223.650 ;
        RECT 106.060 223.615 125.010 223.915 ;
        RECT 103.350 223.015 120.980 223.315 ;
        RECT 100.590 222.415 116.950 222.715 ;
        RECT 97.830 221.815 112.920 222.115 ;
        RECT 95.070 221.215 108.890 221.515 ;
        RECT 92.260 220.510 93.060 220.910 ;
        RECT 1.000 218.590 12.150 220.190 ;
        RECT 106.340 217.515 107.940 219.915 ;
        RECT 6.200 211.890 7.800 215.090 ;
        RECT 9.570 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 9.920 188.640 10.720 211.890 ;
        RECT 15.720 198.970 38.920 209.370 ;
        RECT 9.520 187.840 11.120 188.640 ;
        RECT 15.720 186.970 38.920 197.370 ;
        RECT 44.120 188.440 44.920 211.890 ;
        RECT 6.200 180.050 7.800 183.250 ;
        RECT 9.520 182.990 11.120 183.790 ;
        RECT 3.600 176.050 7.510 179.250 ;
        RECT 9.920 163.040 10.720 182.990 ;
        RECT 15.720 174.970 38.920 185.370 ;
        RECT 45.870 181.190 46.670 210.555 ;
        RECT 106.415 210.540 108.015 213.740 ;
        RECT 47.470 182.790 48.270 204.590 ;
        RECT 108.590 202.625 108.890 221.215 ;
        RECT 109.240 207.925 109.640 219.305 ;
        RECT 110.530 217.705 110.930 219.305 ;
        RECT 110.530 209.640 110.930 211.240 ;
        RECT 111.820 207.925 112.220 219.305 ;
        RECT 109.240 207.525 110.490 207.925 ;
        RECT 108.540 201.825 108.940 202.625 ;
        RECT 63.550 200.610 98.400 200.615 ;
        RECT 63.550 199.815 106.330 200.610 ;
        RECT 98.400 199.810 106.330 199.815 ;
        RECT 68.970 196.830 100.300 197.630 ;
        RECT 74.545 193.735 98.000 194.535 ;
        RECT 66.295 190.655 95.650 191.455 ;
        RECT 52.860 188.465 53.660 190.065 ;
        RECT 55.320 184.940 56.920 186.540 ;
        RECT 47.470 181.990 54.670 182.790 ;
        RECT 45.870 180.390 53.020 181.190 ;
        RECT 9.520 162.240 11.120 163.040 ;
        RECT 15.720 162.970 38.920 173.370 ;
        RECT 52.220 170.440 53.020 180.390 ;
        RECT 53.870 175.290 54.670 181.990 ;
        RECT 53.870 164.840 54.670 174.240 ;
        RECT 55.720 166.640 56.520 184.940 ;
        RECT 57.020 177.390 57.820 178.990 ;
        RECT 61.980 174.370 90.220 175.170 ;
        RECT 57.020 168.290 57.820 169.890 ;
        RECT 55.320 165.840 56.920 166.640 ;
        RECT 53.470 164.040 55.070 164.840 ;
        RECT 9.920 153.790 10.720 162.240 ;
        RECT 9.520 152.990 11.120 153.790 ;
        RECT 9.920 152.915 10.720 152.990 ;
        RECT 15.720 150.970 38.920 161.370 ;
        RECT 51.570 160.190 53.170 160.990 ;
        RECT 51.970 155.790 52.770 160.190 ;
        RECT 51.570 154.990 53.170 155.790 ;
        RECT 41.830 149.410 46.630 150.210 ;
        RECT 51.970 148.290 52.770 154.990 ;
        RECT 53.870 151.990 54.670 164.040 ;
        RECT 53.470 151.190 55.070 151.990 ;
        RECT 55.720 150.240 56.520 165.840 ;
        RECT 54.920 149.440 56.520 150.240 ;
        RECT 51.580 145.090 53.180 148.290 ;
        RECT 61.980 143.690 62.780 174.370 ;
        RECT 3.600 132.225 7.510 135.425 ;
        RECT 9.095 134.635 18.955 143.035 ;
        RECT 20.350 141.375 20.750 142.975 ;
        RECT 28.140 142.890 62.780 143.690 ;
        RECT 13.385 132.330 14.185 133.130 ;
        RECT 20.650 131.410 21.050 138.770 ;
        RECT 61.980 135.095 62.780 142.890 ;
        RECT 70.165 172.130 84.650 172.930 ;
        RECT 22.615 133.320 23.415 134.120 ;
        RECT 16.805 128.710 17.605 129.110 ;
        RECT 6.200 124.285 7.800 127.485 ;
        RECT 12.915 45.565 14.515 119.215 ;
        RECT 16.165 56.765 17.765 121.615 ;
        RECT 21.615 95.165 22.415 132.545 ;
        RECT 27.065 95.165 27.865 130.795 ;
        RECT 70.165 128.125 70.965 172.130 ;
        RECT 74.940 154.795 86.100 155.595 ;
        RECT 71.585 145.090 73.185 148.290 ;
        RECT 74.940 145.235 75.740 154.795 ;
        RECT 94.850 150.520 95.650 190.655 ;
        RECT 80.010 149.520 95.650 150.520 ;
        RECT 74.940 144.435 86.100 145.235 ;
        RECT 63.315 103.770 64.915 123.715 ;
        RECT 65.865 110.280 67.465 127.485 ;
        RECT 75.510 123.715 77.110 135.155 ;
        RECT 80.125 133.320 80.925 144.435 ;
        RECT 94.850 131.745 95.650 149.520 ;
        RECT 97.200 137.420 98.000 193.735 ;
        RECT 99.500 129.995 100.300 196.830 ;
        RECT 102.950 168.255 103.750 186.540 ;
        RECT 105.530 170.890 106.330 199.810 ;
        RECT 109.240 198.885 109.640 205.545 ;
        RECT 110.090 197.895 110.490 207.525 ;
        RECT 109.240 197.495 110.490 197.895 ;
        RECT 110.970 207.525 112.220 207.925 ;
        RECT 110.970 197.895 111.370 207.525 ;
        RECT 111.820 198.885 112.220 206.755 ;
        RECT 112.620 202.625 112.920 221.815 ;
        RECT 113.270 207.925 113.670 219.305 ;
        RECT 114.560 217.705 114.960 219.305 ;
        RECT 114.560 209.640 114.960 211.240 ;
        RECT 115.850 207.925 116.250 219.305 ;
        RECT 113.270 207.525 114.520 207.925 ;
        RECT 112.570 201.825 112.970 202.625 ;
        RECT 113.270 198.885 113.670 205.545 ;
        RECT 114.120 197.895 114.520 207.525 ;
        RECT 110.970 197.495 112.220 197.895 ;
        RECT 109.240 183.970 109.640 197.495 ;
        RECT 111.820 191.285 112.220 197.495 ;
        RECT 113.270 197.495 114.520 197.895 ;
        RECT 115.000 207.525 116.250 207.925 ;
        RECT 115.000 197.895 115.400 207.525 ;
        RECT 115.850 198.885 116.250 206.755 ;
        RECT 116.650 202.625 116.950 222.415 ;
        RECT 117.300 207.925 117.700 219.305 ;
        RECT 118.590 217.705 118.990 219.305 ;
        RECT 118.590 209.640 118.990 211.240 ;
        RECT 119.880 207.925 120.280 219.305 ;
        RECT 117.300 207.525 118.550 207.925 ;
        RECT 116.600 201.825 117.000 202.625 ;
        RECT 117.300 198.885 117.700 205.545 ;
        RECT 118.150 197.895 118.550 207.525 ;
        RECT 115.000 197.495 116.250 197.895 ;
        RECT 110.530 187.540 110.930 189.140 ;
        RECT 113.270 183.990 113.670 197.495 ;
        RECT 115.850 191.285 116.250 197.495 ;
        RECT 117.300 197.495 118.550 197.895 ;
        RECT 119.030 207.525 120.280 207.925 ;
        RECT 119.030 197.895 119.430 207.525 ;
        RECT 119.880 198.885 120.280 206.755 ;
        RECT 120.680 202.625 120.980 223.015 ;
        RECT 121.330 207.925 121.730 219.305 ;
        RECT 122.620 217.705 123.020 219.305 ;
        RECT 122.620 209.640 123.020 211.240 ;
        RECT 123.910 207.925 124.310 219.305 ;
        RECT 121.330 207.525 122.580 207.925 ;
        RECT 120.630 201.825 121.030 202.625 ;
        RECT 121.330 198.885 121.730 205.545 ;
        RECT 122.180 197.895 122.580 207.525 ;
        RECT 119.030 197.495 120.280 197.895 ;
        RECT 114.560 187.540 114.960 189.140 ;
        RECT 111.685 183.590 113.670 183.990 ;
        RECT 105.530 168.255 106.730 170.890 ;
        RECT 107.380 168.490 107.780 170.890 ;
        RECT 103.350 152.765 103.750 160.495 ;
        RECT 103.350 143.435 103.750 145.835 ;
        RECT 104.640 140.165 105.040 167.190 ;
        RECT 105.385 157.365 105.785 158.165 ;
        RECT 106.330 145.835 106.730 168.255 ;
        RECT 107.380 152.765 107.780 160.495 ;
        RECT 108.670 147.135 109.070 178.990 ;
        RECT 109.960 168.490 110.760 170.890 ;
        RECT 109.415 156.165 109.815 156.965 ;
        RECT 110.360 145.835 110.760 168.490 ;
        RECT 111.685 157.765 112.085 183.590 ;
        RECT 117.300 182.580 117.700 197.495 ;
        RECT 119.880 191.285 120.280 197.495 ;
        RECT 121.330 197.495 122.580 197.895 ;
        RECT 123.060 207.525 124.310 207.925 ;
        RECT 123.060 197.895 123.460 207.525 ;
        RECT 123.910 198.885 124.310 206.755 ;
        RECT 124.710 202.625 125.010 223.615 ;
        RECT 125.360 207.925 125.760 219.305 ;
        RECT 126.650 217.705 127.050 219.305 ;
        RECT 126.650 209.640 127.050 211.240 ;
        RECT 127.940 207.925 128.340 219.305 ;
        RECT 125.360 207.525 126.610 207.925 ;
        RECT 124.660 201.825 125.060 202.625 ;
        RECT 125.360 198.885 125.760 205.545 ;
        RECT 126.210 197.895 126.610 207.525 ;
        RECT 123.060 197.495 124.310 197.895 ;
        RECT 118.590 187.540 118.990 189.140 ;
        RECT 113.085 182.180 117.700 182.580 ;
        RECT 113.085 156.165 113.485 182.180 ;
        RECT 121.330 181.545 121.730 197.495 ;
        RECT 123.910 191.285 124.310 197.495 ;
        RECT 125.360 197.495 126.610 197.895 ;
        RECT 127.090 207.525 128.340 207.925 ;
        RECT 127.090 197.895 127.490 207.525 ;
        RECT 127.940 198.885 128.340 206.755 ;
        RECT 128.740 202.625 129.040 224.215 ;
        RECT 132.720 220.715 133.120 221.515 ;
        RECT 136.750 220.715 137.150 221.515 ;
        RECT 140.780 220.715 141.180 221.515 ;
        RECT 144.810 220.715 145.210 221.515 ;
        RECT 148.840 220.715 149.240 221.515 ;
        RECT 129.390 207.925 129.790 219.305 ;
        RECT 130.680 217.705 131.080 219.305 ;
        RECT 130.680 209.640 131.080 211.240 ;
        RECT 131.970 207.925 132.370 219.305 ;
        RECT 129.390 207.525 130.640 207.925 ;
        RECT 128.690 201.825 129.090 202.625 ;
        RECT 129.390 198.885 129.790 205.545 ;
        RECT 130.240 197.895 130.640 207.525 ;
        RECT 127.090 197.495 128.340 197.895 ;
        RECT 122.620 187.540 123.020 189.140 ;
        RECT 116.415 181.145 121.730 181.545 ;
        RECT 116.415 176.215 116.815 181.145 ;
        RECT 125.360 180.565 125.760 197.495 ;
        RECT 127.940 191.285 128.340 197.495 ;
        RECT 129.390 197.495 130.640 197.895 ;
        RECT 131.120 207.525 132.370 207.925 ;
        RECT 131.120 197.895 131.520 207.525 ;
        RECT 131.970 198.885 132.370 206.755 ;
        RECT 132.770 202.625 133.070 220.715 ;
        RECT 133.420 207.925 133.820 219.305 ;
        RECT 134.710 217.705 135.110 219.305 ;
        RECT 134.710 209.640 135.110 211.240 ;
        RECT 136.000 207.925 136.400 219.305 ;
        RECT 133.420 207.525 134.670 207.925 ;
        RECT 132.720 201.825 133.120 202.625 ;
        RECT 133.420 198.885 133.820 205.545 ;
        RECT 134.270 197.895 134.670 207.525 ;
        RECT 131.120 197.495 132.370 197.895 ;
        RECT 126.650 187.540 127.050 189.140 ;
        RECT 121.035 180.165 125.760 180.565 ;
        RECT 121.035 176.215 121.435 180.165 ;
        RECT 129.390 179.490 129.790 197.495 ;
        RECT 131.970 191.285 132.370 197.495 ;
        RECT 133.420 197.495 134.670 197.895 ;
        RECT 135.150 207.525 136.400 207.925 ;
        RECT 135.150 197.895 135.550 207.525 ;
        RECT 136.000 198.885 136.400 206.755 ;
        RECT 136.800 202.625 137.100 220.715 ;
        RECT 137.450 207.925 137.850 219.305 ;
        RECT 138.740 217.705 139.140 219.305 ;
        RECT 138.740 209.640 139.140 211.240 ;
        RECT 140.030 207.925 140.430 219.305 ;
        RECT 137.450 207.525 138.700 207.925 ;
        RECT 136.750 201.825 137.150 202.625 ;
        RECT 137.450 198.885 137.850 205.545 ;
        RECT 138.300 197.895 138.700 207.525 ;
        RECT 135.150 197.495 136.400 197.895 ;
        RECT 130.680 187.540 131.080 189.140 ;
        RECT 125.660 179.090 129.790 179.490 ;
        RECT 125.660 176.215 126.060 179.090 ;
        RECT 133.420 178.920 133.820 197.495 ;
        RECT 136.000 191.285 136.400 197.495 ;
        RECT 137.450 197.495 138.700 197.895 ;
        RECT 139.180 207.525 140.430 207.925 ;
        RECT 139.180 197.895 139.580 207.525 ;
        RECT 140.030 198.885 140.430 206.755 ;
        RECT 140.830 202.625 141.130 220.715 ;
        RECT 141.480 207.925 141.880 219.305 ;
        RECT 142.770 217.705 143.170 219.305 ;
        RECT 142.770 209.640 143.170 211.240 ;
        RECT 144.060 207.925 144.460 219.305 ;
        RECT 141.480 207.525 142.730 207.925 ;
        RECT 140.780 201.825 141.180 202.625 ;
        RECT 141.480 198.885 141.880 205.545 ;
        RECT 142.330 197.895 142.730 207.525 ;
        RECT 139.180 197.495 140.430 197.895 ;
        RECT 134.710 187.540 135.110 189.140 ;
        RECT 137.450 178.920 137.850 197.495 ;
        RECT 140.030 191.285 140.430 197.495 ;
        RECT 141.480 197.495 142.730 197.895 ;
        RECT 143.210 207.525 144.460 207.925 ;
        RECT 143.210 197.895 143.610 207.525 ;
        RECT 144.060 198.885 144.460 206.755 ;
        RECT 144.860 202.625 145.160 220.715 ;
        RECT 145.510 207.925 145.910 219.305 ;
        RECT 146.800 217.705 147.200 219.305 ;
        RECT 146.800 209.640 147.200 211.240 ;
        RECT 148.090 207.925 148.490 219.305 ;
        RECT 145.510 207.525 146.760 207.925 ;
        RECT 144.810 201.825 145.210 202.625 ;
        RECT 145.510 198.885 145.910 205.545 ;
        RECT 146.360 197.895 146.760 207.525 ;
        RECT 143.210 197.495 144.460 197.895 ;
        RECT 138.740 187.540 139.140 189.140 ;
        RECT 141.480 178.920 141.880 197.495 ;
        RECT 144.060 191.285 144.460 197.495 ;
        RECT 145.510 197.495 146.760 197.895 ;
        RECT 147.240 207.525 148.490 207.925 ;
        RECT 147.240 197.895 147.640 207.525 ;
        RECT 148.090 198.885 148.490 206.755 ;
        RECT 148.890 202.625 149.190 220.715 ;
        RECT 162.100 220.260 162.500 220.910 ;
        RECT 163.100 220.860 163.500 221.510 ;
        RECT 164.100 221.460 164.500 222.110 ;
        RECT 164.100 221.160 250.220 221.460 ;
        RECT 163.100 220.560 249.370 220.860 ;
        RECT 162.100 219.960 248.285 220.260 ;
        RECT 149.540 207.925 149.940 219.305 ;
        RECT 150.830 217.705 151.230 219.305 ;
        RECT 150.830 209.640 151.230 211.240 ;
        RECT 152.120 207.925 152.520 219.305 ;
        RECT 246.615 217.650 247.015 218.450 ;
        RECT 149.540 207.525 150.790 207.925 ;
        RECT 148.840 201.825 149.240 202.625 ;
        RECT 149.540 198.885 149.940 205.545 ;
        RECT 150.390 197.895 150.790 207.525 ;
        RECT 147.240 197.495 148.490 197.895 ;
        RECT 142.770 187.540 143.170 189.140 ;
        RECT 145.510 178.920 145.910 197.495 ;
        RECT 148.090 191.285 148.490 197.495 ;
        RECT 149.540 197.495 150.790 197.895 ;
        RECT 151.270 207.525 152.520 207.925 ;
        RECT 151.270 197.895 151.670 207.525 ;
        RECT 152.120 198.885 152.520 206.755 ;
        RECT 180.680 201.325 182.260 201.655 ;
        RECT 183.980 198.605 185.560 198.935 ;
        RECT 162.390 197.900 164.390 198.050 ;
        RECT 166.595 197.900 166.925 197.915 ;
        RECT 151.270 197.495 152.520 197.895 ;
        RECT 146.800 187.540 147.200 189.140 ;
        RECT 149.540 178.920 149.940 197.495 ;
        RECT 152.120 191.285 152.520 197.495 ;
        RECT 159.185 197.600 166.925 197.900 ;
        RECT 150.830 187.540 151.230 189.140 ;
        RECT 153.565 184.765 155.165 187.965 ;
        RECT 158.335 187.580 158.735 188.380 ;
        RECT 130.275 178.520 133.820 178.920 ;
        RECT 134.895 178.520 137.850 178.920 ;
        RECT 139.510 178.520 141.880 178.920 ;
        RECT 144.135 178.520 145.910 178.920 ;
        RECT 148.755 178.520 149.940 178.920 ;
        RECT 130.275 176.215 130.675 178.520 ;
        RECT 134.895 176.215 135.295 178.520 ;
        RECT 139.510 176.215 139.910 178.520 ;
        RECT 144.135 176.215 144.535 178.520 ;
        RECT 148.755 176.215 149.155 178.520 ;
        RECT 116.215 175.815 117.015 176.215 ;
        RECT 120.835 175.815 121.635 176.215 ;
        RECT 125.455 175.815 126.255 176.215 ;
        RECT 130.075 175.815 130.875 176.215 ;
        RECT 134.695 175.815 135.495 176.215 ;
        RECT 139.315 175.815 140.115 176.215 ;
        RECT 143.935 175.815 144.735 176.215 ;
        RECT 148.555 175.815 149.355 176.215 ;
        RECT 151.155 175.010 152.755 178.210 ;
        RECT 115.815 173.070 117.415 173.870 ;
        RECT 120.435 173.070 122.035 173.870 ;
        RECT 125.055 173.070 126.655 173.870 ;
        RECT 129.675 173.070 131.275 173.870 ;
        RECT 134.295 173.070 135.895 173.870 ;
        RECT 138.915 173.070 140.515 173.870 ;
        RECT 143.535 173.070 145.135 173.870 ;
        RECT 148.155 173.070 149.755 173.870 ;
        RECT 105.930 143.435 106.730 145.835 ;
        RECT 104.640 139.365 105.440 140.165 ;
        RECT 107.380 136.325 107.780 145.835 ;
        RECT 109.960 143.435 110.760 145.835 ;
        RECT 116.310 144.730 116.910 173.070 ;
        RECT 120.930 147.530 121.530 173.070 ;
        RECT 125.550 148.690 126.150 173.070 ;
        RECT 130.175 149.890 130.775 173.070 ;
        RECT 134.795 160.260 135.395 173.070 ;
        RECT 136.775 161.650 137.575 162.450 ;
        RECT 134.695 159.460 135.495 160.260 ;
        RECT 133.275 152.100 134.875 152.200 ;
        RECT 136.875 152.100 137.475 161.650 ;
        RECT 133.275 151.500 137.475 152.100 ;
        RECT 133.275 151.400 134.875 151.500 ;
        RECT 133.275 150.930 134.875 151.030 ;
        RECT 139.410 150.930 140.010 173.070 ;
        RECT 144.035 162.450 144.635 173.070 ;
        RECT 143.935 161.650 144.735 162.450 ;
        RECT 148.655 161.210 149.255 173.070 ;
        RECT 133.275 150.330 140.010 150.930 ;
        RECT 141.715 160.610 149.255 161.210 ;
        RECT 133.275 150.230 134.875 150.330 ;
        RECT 130.175 149.290 136.695 149.890 ;
        RECT 125.550 148.090 133.635 148.690 ;
        RECT 130.615 147.530 132.215 147.630 ;
        RECT 120.930 146.930 132.215 147.530 ;
        RECT 130.615 146.830 132.215 146.930 ;
        RECT 122.645 144.730 124.245 144.830 ;
        RECT 116.310 144.130 124.245 144.730 ;
        RECT 122.645 144.030 124.245 144.130 ;
        RECT 133.035 144.520 133.635 148.090 ;
        RECT 136.095 148.010 136.695 149.290 ;
        RECT 138.525 148.010 140.125 148.110 ;
        RECT 136.095 147.410 140.125 148.010 ;
        RECT 138.525 147.310 140.125 147.410 ;
        RECT 138.525 144.520 140.125 144.620 ;
        RECT 133.035 143.920 140.125 144.520 ;
        RECT 141.715 144.040 142.315 160.610 ;
        RECT 145.525 159.460 146.325 160.260 ;
        RECT 138.525 143.820 140.125 143.920 ;
        RECT 109.960 138.220 110.360 143.435 ;
        RECT 141.215 143.240 142.815 144.040 ;
        RECT 141.215 142.690 142.815 142.790 ;
        RECT 145.625 142.690 146.225 159.460 ;
        RECT 141.215 142.090 146.225 142.690 ;
        RECT 141.215 141.990 142.815 142.090 ;
        RECT 109.560 137.420 110.760 138.220 ;
        RECT 107.380 135.525 108.180 136.325 ;
        RECT 72.765 103.865 74.365 122.215 ;
        RECT 75.510 114.215 77.115 123.715 ;
        RECT 75.515 100.215 77.115 114.215 ;
        RECT 21.215 51.675 22.815 95.165 ;
        RECT 26.665 61.465 28.265 95.165 ;
        RECT 97.165 93.265 98.765 119.215 ;
        RECT 100.515 117.715 101.315 128.925 ;
        RECT 100.115 96.415 101.715 117.715 ;
        RECT 103.315 111.365 104.915 123.165 ;
        RECT 116.915 121.965 118.515 122.765 ;
        RECT 105.965 103.965 107.565 120.665 ;
        RECT 109.865 108.365 111.465 119.215 ;
        RECT 117.115 108.365 118.715 118.265 ;
        RECT 121.565 113.015 123.165 127.485 ;
        RECT 116.965 104.015 118.565 104.815 ;
        RECT 42.740 71.190 53.140 83.050 ;
        RECT 55.740 71.190 66.140 83.050 ;
        RECT 68.740 71.190 79.140 83.050 ;
        RECT 81.740 71.190 92.140 83.050 ;
        RECT 94.740 71.190 105.140 83.050 ;
        RECT 42.740 57.830 53.140 69.690 ;
        RECT 55.740 57.830 66.140 69.690 ;
        RECT 68.740 57.830 79.140 69.690 ;
        RECT 81.740 57.830 92.140 69.690 ;
        RECT 94.740 57.830 105.140 69.690 ;
        RECT 6.200 41.635 7.800 44.835 ;
        RECT 3.600 36.430 8.665 39.630 ;
        RECT 3.600 5.690 8.665 8.890 ;
        RECT 14.965 5.690 16.565 34.940 ;
        RECT 65.765 15.915 67.365 44.215 ;
        RECT 68.865 11.965 70.465 41.615 ;
        RECT 72.095 9.665 73.695 38.865 ;
        RECT 80.745 9.665 82.345 37.635 ;
        RECT 84.015 22.315 85.615 41.615 ;
        RECT 87.165 26.815 88.765 44.215 ;
        RECT 90.715 19.315 92.315 47.165 ;
        RECT 116.115 42.615 117.715 90.815 ;
        RECT 119.215 40.015 120.815 84.315 ;
        RECT 123.215 23.815 124.815 94.865 ;
        RECT 126.165 25.365 127.765 98.015 ;
        RECT 128.965 5.690 130.565 8.890 ;
        RECT 2.705 1.285 98.380 2.085 ;
        RECT 131.665 1.800 132.465 136.325 ;
        RECT 133.265 111.795 134.065 130.795 ;
        RECT 134.865 110.315 135.665 132.545 ;
        RECT 136.465 114.770 137.265 134.120 ;
        RECT 137.945 133.410 138.745 133.810 ;
        RECT 137.945 131.410 138.345 133.410 ;
        RECT 139.120 131.390 139.520 132.990 ;
        RECT 141.700 131.390 142.100 132.990 ;
        RECT 139.120 125.690 139.520 127.290 ;
        RECT 139.970 125.690 142.100 127.290 ;
        RECT 142.760 122.490 145.960 124.090 ;
        RECT 133.525 109.515 138.400 110.315 ;
        RECT 136.295 108.925 138.400 109.515 ;
        RECT 136.295 94.305 138.400 94.895 ;
        RECT 136.495 29.375 138.195 94.305 ;
        RECT 139.355 30.545 141.055 114.150 ;
        RECT 141.900 110.315 142.700 117.170 ;
        RECT 138.950 29.955 141.055 30.545 ;
        RECT 136.295 28.785 138.400 29.375 ;
        RECT 141.495 20.015 143.195 110.315 ;
        RECT 143.640 32.885 145.340 114.150 ;
        RECT 146.950 110.315 147.750 138.220 ;
        RECT 149.945 116.370 150.745 170.845 ;
        RECT 146.490 104.255 148.190 110.315 ;
        RECT 146.290 103.665 148.395 104.255 ;
        RECT 143.640 32.295 145.745 32.885 ;
        RECT 141.295 19.425 143.400 20.015 ;
        RECT 151.560 1.800 152.360 140.165 ;
        RECT 153.945 129.145 154.345 184.370 ;
        RECT 157.560 178.060 157.960 178.860 ;
        RECT 157.560 28.035 157.860 178.060 ;
        RECT 158.335 60.675 158.635 187.580 ;
        RECT 159.185 93.465 159.485 197.600 ;
        RECT 162.390 197.450 164.390 197.600 ;
        RECT 166.595 197.585 166.925 197.600 ;
        RECT 180.680 195.885 182.260 196.215 ;
        RECT 183.980 193.165 185.560 193.495 ;
        RECT 167.515 193.140 167.845 193.155 ;
        RECT 181.775 193.140 182.105 193.155 ;
        RECT 167.515 192.840 182.105 193.140 ;
        RECT 167.515 192.825 167.845 192.840 ;
        RECT 181.775 192.825 182.105 192.840 ;
        RECT 174.415 192.460 174.745 192.475 ;
        RECT 184.075 192.460 184.405 192.475 ;
        RECT 174.415 192.160 184.405 192.460 ;
        RECT 174.415 192.145 174.745 192.160 ;
        RECT 184.075 192.145 184.405 192.160 ;
        RECT 179.015 191.780 179.345 191.795 ;
        RECT 193.735 191.780 194.065 191.795 ;
        RECT 179.015 191.480 194.065 191.780 ;
        RECT 179.015 191.465 179.345 191.480 ;
        RECT 193.735 191.465 194.065 191.480 ;
        RECT 180.680 190.445 182.260 190.775 ;
        RECT 177.380 189.740 177.760 189.750 ;
        RECT 196.495 189.740 196.825 189.755 ;
        RECT 177.380 189.440 196.825 189.740 ;
        RECT 177.380 189.430 177.760 189.440 ;
        RECT 196.495 189.425 196.825 189.440 ;
        RECT 179.015 189.060 179.345 189.075 ;
        RECT 184.995 189.060 185.325 189.075 ;
        RECT 179.015 188.760 185.325 189.060 ;
        RECT 179.015 188.745 179.345 188.760 ;
        RECT 184.995 188.745 185.325 188.760 ;
        RECT 162.390 188.430 164.390 188.530 ;
        RECT 161.590 188.380 164.390 188.430 ;
        RECT 166.595 188.380 166.925 188.395 ;
        RECT 161.590 188.080 166.925 188.380 ;
        RECT 161.590 188.030 164.390 188.080 ;
        RECT 166.595 188.065 166.925 188.080 ;
        RECT 162.390 187.930 164.390 188.030 ;
        RECT 183.980 187.725 185.560 188.055 ;
        RECT 167.975 187.700 168.305 187.715 ;
        RECT 179.935 187.700 180.265 187.715 ;
        RECT 167.975 187.400 180.265 187.700 ;
        RECT 167.975 187.385 168.305 187.400 ;
        RECT 179.935 187.385 180.265 187.400 ;
        RECT 230.535 187.700 230.865 187.715 ;
        RECT 232.835 187.700 233.165 187.715 ;
        RECT 230.535 187.400 233.165 187.700 ;
        RECT 230.535 187.385 230.865 187.400 ;
        RECT 232.835 187.385 233.165 187.400 ;
        RECT 180.395 187.020 180.725 187.035 ;
        RECT 200.175 187.020 200.505 187.035 ;
        RECT 180.395 186.720 200.505 187.020 ;
        RECT 180.395 186.705 180.725 186.720 ;
        RECT 200.175 186.705 200.505 186.720 ;
        RECT 201.095 187.020 201.425 187.035 ;
        RECT 233.755 187.020 234.085 187.035 ;
        RECT 201.095 186.720 234.085 187.020 ;
        RECT 201.095 186.705 201.425 186.720 ;
        RECT 233.755 186.705 234.085 186.720 ;
        RECT 179.220 186.340 179.600 186.350 ;
        RECT 187.295 186.340 187.625 186.355 ;
        RECT 179.220 186.040 187.625 186.340 ;
        RECT 179.220 186.030 179.600 186.040 ;
        RECT 187.295 186.025 187.625 186.040 ;
        RECT 209.835 186.340 210.165 186.355 ;
        RECT 236.515 186.340 236.845 186.355 ;
        RECT 209.835 186.040 236.845 186.340 ;
        RECT 209.835 186.025 210.165 186.040 ;
        RECT 236.515 186.025 236.845 186.040 ;
        RECT 190.055 185.670 190.385 185.675 ;
        RECT 190.055 185.660 190.640 185.670 ;
        RECT 213.055 185.660 213.385 185.675 ;
        RECT 190.055 185.360 190.840 185.660 ;
        RECT 210.540 185.360 213.385 185.660 ;
        RECT 190.055 185.350 190.640 185.360 ;
        RECT 190.055 185.345 190.385 185.350 ;
        RECT 180.680 185.005 182.260 185.335 ;
        RECT 175.540 184.300 175.920 184.310 ;
        RECT 177.175 184.300 177.505 184.315 ;
        RECT 175.540 184.000 177.505 184.300 ;
        RECT 175.540 183.990 175.920 184.000 ;
        RECT 177.175 183.985 177.505 184.000 ;
        RECT 182.900 184.300 183.280 184.310 ;
        RECT 184.995 184.300 185.325 184.315 ;
        RECT 182.900 184.000 185.325 184.300 ;
        RECT 182.900 183.990 183.280 184.000 ;
        RECT 184.995 183.985 185.325 184.000 ;
        RECT 186.835 184.300 187.165 184.315 ;
        RECT 190.975 184.300 191.305 184.315 ;
        RECT 186.835 184.000 191.305 184.300 ;
        RECT 186.835 183.985 187.165 184.000 ;
        RECT 190.975 183.985 191.305 184.000 ;
        RECT 175.795 183.620 176.125 183.635 ;
        RECT 181.315 183.620 181.645 183.635 ;
        RECT 189.595 183.620 189.925 183.635 ;
        RECT 175.795 183.320 189.925 183.620 ;
        RECT 175.795 183.305 176.125 183.320 ;
        RECT 181.315 183.305 181.645 183.320 ;
        RECT 189.595 183.305 189.925 183.320 ;
        RECT 175.795 182.940 176.125 182.955 ;
        RECT 176.715 182.940 177.045 182.955 ;
        RECT 175.795 182.640 177.045 182.940 ;
        RECT 175.795 182.625 176.125 182.640 ;
        RECT 176.715 182.625 177.045 182.640 ;
        RECT 186.835 182.940 187.165 182.955 ;
        RECT 192.355 182.940 192.685 182.955 ;
        RECT 186.835 182.640 192.685 182.940 ;
        RECT 186.835 182.625 187.165 182.640 ;
        RECT 192.355 182.625 192.685 182.640 ;
        RECT 183.980 182.285 185.560 182.615 ;
        RECT 210.540 182.275 210.840 185.360 ;
        RECT 213.055 185.345 213.385 185.360 ;
        RECT 212.340 184.980 212.720 184.990 ;
        RECT 234.215 184.980 234.545 184.995 ;
        RECT 212.340 184.680 234.545 184.980 ;
        RECT 212.340 184.670 212.720 184.680 ;
        RECT 234.215 184.665 234.545 184.680 ;
        RECT 223.635 183.620 223.965 183.635 ;
        RECT 224.555 183.620 224.885 183.635 ;
        RECT 223.635 183.320 224.885 183.620 ;
        RECT 223.635 183.305 223.965 183.320 ;
        RECT 224.555 183.305 224.885 183.320 ;
        RECT 227.315 183.620 227.645 183.635 ;
        RECT 230.075 183.620 230.405 183.635 ;
        RECT 227.315 183.320 230.405 183.620 ;
        RECT 227.315 183.305 227.645 183.320 ;
        RECT 230.075 183.305 230.405 183.320 ;
        RECT 211.675 182.940 212.005 182.955 ;
        RECT 232.375 182.940 232.705 182.955 ;
        RECT 211.675 182.640 232.705 182.940 ;
        RECT 211.675 182.625 212.005 182.640 ;
        RECT 232.375 182.625 232.705 182.640 ;
        RECT 186.375 182.260 186.705 182.275 ;
        RECT 200.175 182.260 200.505 182.275 ;
        RECT 186.375 181.960 200.505 182.260 ;
        RECT 210.540 181.960 211.085 182.275 ;
        RECT 186.375 181.945 186.705 181.960 ;
        RECT 200.175 181.945 200.505 181.960 ;
        RECT 210.755 181.945 211.085 181.960 ;
        RECT 211.675 182.260 212.005 182.275 ;
        RECT 232.835 182.260 233.165 182.275 ;
        RECT 211.675 181.960 233.165 182.260 ;
        RECT 211.675 181.945 212.005 181.960 ;
        RECT 232.835 181.945 233.165 181.960 ;
        RECT 169.355 181.580 169.685 181.595 ;
        RECT 175.795 181.580 176.125 181.595 ;
        RECT 169.355 181.280 176.125 181.580 ;
        RECT 169.355 181.265 169.685 181.280 ;
        RECT 175.795 181.265 176.125 181.280 ;
        RECT 182.235 181.580 182.565 181.595 ;
        RECT 186.835 181.580 187.165 181.595 ;
        RECT 182.235 181.280 187.165 181.580 ;
        RECT 182.235 181.265 182.565 181.280 ;
        RECT 186.835 181.265 187.165 181.280 ;
        RECT 190.515 181.580 190.845 181.595 ;
        RECT 198.795 181.580 199.125 181.595 ;
        RECT 190.515 181.280 199.125 181.580 ;
        RECT 190.515 181.265 190.845 181.280 ;
        RECT 198.795 181.265 199.125 181.280 ;
        RECT 210.295 181.580 210.625 181.595 ;
        RECT 227.775 181.580 228.105 181.595 ;
        RECT 234.675 181.580 235.005 181.595 ;
        RECT 210.295 181.280 227.400 181.580 ;
        RECT 210.295 181.265 210.625 181.280 ;
        RECT 172.115 180.900 172.445 180.915 ;
        RECT 216.275 180.900 216.605 180.915 ;
        RECT 172.115 180.600 216.605 180.900 ;
        RECT 227.100 180.900 227.400 181.280 ;
        RECT 227.775 181.280 235.005 181.580 ;
        RECT 227.775 181.265 228.105 181.280 ;
        RECT 234.675 181.265 235.005 181.280 ;
        RECT 227.775 180.900 228.105 180.915 ;
        RECT 227.100 180.600 228.105 180.900 ;
        RECT 172.115 180.585 172.445 180.600 ;
        RECT 216.275 180.585 216.605 180.600 ;
        RECT 227.775 180.585 228.105 180.600 ;
        RECT 168.895 180.220 169.225 180.235 ;
        RECT 179.015 180.220 179.345 180.235 ;
        RECT 168.895 179.920 179.345 180.220 ;
        RECT 168.895 179.905 169.225 179.920 ;
        RECT 179.015 179.905 179.345 179.920 ;
        RECT 182.900 180.220 183.280 180.230 ;
        RECT 183.615 180.220 183.945 180.235 ;
        RECT 182.900 179.920 183.945 180.220 ;
        RECT 182.900 179.910 183.280 179.920 ;
        RECT 183.615 179.905 183.945 179.920 ;
        RECT 184.535 180.220 184.865 180.235 ;
        RECT 196.035 180.220 196.365 180.235 ;
        RECT 184.535 179.920 196.365 180.220 ;
        RECT 184.535 179.905 184.865 179.920 ;
        RECT 196.035 179.905 196.365 179.920 ;
        RECT 213.975 180.220 214.305 180.235 ;
        RECT 217.195 180.220 217.525 180.235 ;
        RECT 213.975 179.920 217.525 180.220 ;
        RECT 213.975 179.905 214.305 179.920 ;
        RECT 217.195 179.905 217.525 179.920 ;
        RECT 221.795 180.220 222.125 180.235 ;
        RECT 235.595 180.220 235.925 180.235 ;
        RECT 221.795 179.920 235.925 180.220 ;
        RECT 221.795 179.905 222.125 179.920 ;
        RECT 235.595 179.905 235.925 179.920 ;
        RECT 180.680 179.565 182.260 179.895 ;
        RECT 175.335 179.550 175.665 179.555 ;
        RECT 177.635 179.550 177.965 179.555 ;
        RECT 175.335 179.540 175.920 179.550 ;
        RECT 175.110 179.240 175.920 179.540 ;
        RECT 175.335 179.230 175.920 179.240 ;
        RECT 177.380 179.540 177.965 179.550 ;
        RECT 185.455 179.540 185.785 179.555 ;
        RECT 193.735 179.540 194.065 179.555 ;
        RECT 177.380 179.240 178.190 179.540 ;
        RECT 185.455 179.240 194.065 179.540 ;
        RECT 177.380 179.230 177.965 179.240 ;
        RECT 175.335 179.225 175.665 179.230 ;
        RECT 177.635 179.225 177.965 179.230 ;
        RECT 185.455 179.225 185.785 179.240 ;
        RECT 193.735 179.225 194.065 179.240 ;
        RECT 212.135 179.550 212.465 179.555 ;
        RECT 212.135 179.540 212.720 179.550 ;
        RECT 214.435 179.540 214.765 179.555 ;
        RECT 217.655 179.540 217.985 179.555 ;
        RECT 212.135 179.240 212.920 179.540 ;
        RECT 214.435 179.240 217.985 179.540 ;
        RECT 212.135 179.230 212.720 179.240 ;
        RECT 212.135 179.225 212.465 179.230 ;
        RECT 214.435 179.225 214.765 179.240 ;
        RECT 217.655 179.225 217.985 179.240 ;
        RECT 219.035 179.540 219.365 179.555 ;
        RECT 231.455 179.540 231.785 179.555 ;
        RECT 219.035 179.240 231.785 179.540 ;
        RECT 219.035 179.225 219.365 179.240 ;
        RECT 231.455 179.225 231.785 179.240 ;
        RECT 162.390 178.910 164.390 179.010 ;
        RECT 161.590 178.860 164.390 178.910 ;
        RECT 167.055 178.860 167.385 178.875 ;
        RECT 161.590 178.560 167.385 178.860 ;
        RECT 161.590 178.510 164.390 178.560 ;
        RECT 167.055 178.545 167.385 178.560 ;
        RECT 169.355 178.860 169.685 178.875 ;
        RECT 178.555 178.860 178.885 178.875 ;
        RECT 179.220 178.860 179.600 178.870 ;
        RECT 169.355 178.560 176.340 178.860 ;
        RECT 169.355 178.545 169.685 178.560 ;
        RECT 162.390 178.410 164.390 178.510 ;
        RECT 176.040 178.180 176.340 178.560 ;
        RECT 178.555 178.560 179.600 178.860 ;
        RECT 178.555 178.545 178.885 178.560 ;
        RECT 179.220 178.550 179.600 178.560 ;
        RECT 181.315 178.860 181.645 178.875 ;
        RECT 192.355 178.860 192.685 178.875 ;
        RECT 181.315 178.560 192.685 178.860 ;
        RECT 181.315 178.545 181.645 178.560 ;
        RECT 192.355 178.545 192.685 178.560 ;
        RECT 202.935 178.860 203.265 178.875 ;
        RECT 226.395 178.860 226.725 178.875 ;
        RECT 232.835 178.860 233.165 178.875 ;
        RECT 202.935 178.560 226.725 178.860 ;
        RECT 202.935 178.545 203.265 178.560 ;
        RECT 226.395 178.545 226.725 178.560 ;
        RECT 228.940 178.560 233.165 178.860 ;
        RECT 201.095 178.180 201.425 178.195 ;
        RECT 176.040 177.880 201.425 178.180 ;
        RECT 201.095 177.865 201.425 177.880 ;
        RECT 210.295 178.180 210.625 178.195 ;
        RECT 213.055 178.180 213.385 178.195 ;
        RECT 223.175 178.180 223.505 178.195 ;
        RECT 225.935 178.180 226.265 178.195 ;
        RECT 228.940 178.180 229.240 178.560 ;
        RECT 232.835 178.545 233.165 178.560 ;
        RECT 210.295 177.880 229.240 178.180 ;
        RECT 230.075 178.180 230.405 178.195 ;
        RECT 236.055 178.180 236.385 178.195 ;
        RECT 230.075 177.880 236.385 178.180 ;
        RECT 210.295 177.865 210.625 177.880 ;
        RECT 213.055 177.865 213.385 177.880 ;
        RECT 223.175 177.865 223.505 177.880 ;
        RECT 225.935 177.865 226.265 177.880 ;
        RECT 230.075 177.865 230.405 177.880 ;
        RECT 236.055 177.865 236.385 177.880 ;
        RECT 189.595 177.500 189.925 177.515 ;
        RECT 190.260 177.500 190.640 177.510 ;
        RECT 189.595 177.200 190.640 177.500 ;
        RECT 189.595 177.185 189.925 177.200 ;
        RECT 190.260 177.190 190.640 177.200 ;
        RECT 190.975 177.500 191.305 177.515 ;
        RECT 197.875 177.500 198.205 177.515 ;
        RECT 190.975 177.200 198.205 177.500 ;
        RECT 190.975 177.185 191.305 177.200 ;
        RECT 197.875 177.185 198.205 177.200 ;
        RECT 215.355 177.500 215.685 177.515 ;
        RECT 218.575 177.500 218.905 177.515 ;
        RECT 227.775 177.500 228.105 177.515 ;
        RECT 215.355 177.200 218.905 177.500 ;
        RECT 215.355 177.185 215.685 177.200 ;
        RECT 218.575 177.185 218.905 177.200 ;
        RECT 226.180 177.200 228.105 177.500 ;
        RECT 183.980 176.845 185.560 177.175 ;
        RECT 168.435 176.820 168.765 176.835 ;
        RECT 181.315 176.820 181.645 176.835 ;
        RECT 168.435 176.520 181.645 176.820 ;
        RECT 168.435 176.505 168.765 176.520 ;
        RECT 181.315 176.505 181.645 176.520 ;
        RECT 182.695 176.820 183.025 176.835 ;
        RECT 225.475 176.820 225.805 176.835 ;
        RECT 226.180 176.820 226.480 177.200 ;
        RECT 227.775 177.185 228.105 177.200 ;
        RECT 182.695 176.505 183.240 176.820 ;
        RECT 225.475 176.520 226.480 176.820 ;
        RECT 227.315 176.820 227.645 176.835 ;
        RECT 233.295 176.820 233.625 176.835 ;
        RECT 227.315 176.520 233.625 176.820 ;
        RECT 225.475 176.505 225.805 176.520 ;
        RECT 227.315 176.505 227.645 176.520 ;
        RECT 233.295 176.505 233.625 176.520 ;
        RECT 182.940 176.140 183.240 176.505 ;
        RECT 190.975 176.140 191.305 176.155 ;
        RECT 182.940 175.840 191.305 176.140 ;
        RECT 190.975 175.825 191.305 175.840 ;
        RECT 225.015 176.140 225.345 176.155 ;
        RECT 234.215 176.140 234.545 176.155 ;
        RECT 225.015 175.840 234.545 176.140 ;
        RECT 225.015 175.825 225.345 175.840 ;
        RECT 234.215 175.825 234.545 175.840 ;
        RECT 246.665 152.705 246.965 217.650 ;
        RECT 247.985 153.875 248.285 219.960 ;
        RECT 249.070 154.925 249.370 220.560 ;
        RECT 249.920 155.950 250.220 221.160 ;
        RECT 250.925 157.080 251.225 224.750 ;
        RECT 251.860 158.175 252.160 225.410 ;
        RECT 251.860 157.875 318.785 158.175 ;
        RECT 250.925 156.780 317.675 157.080 ;
        RECT 249.920 155.650 316.845 155.950 ;
        RECT 249.070 154.625 316.145 154.925 ;
        RECT 247.985 153.575 315.370 153.875 ;
        RECT 246.665 152.405 314.635 152.705 ;
        RECT 180.925 106.260 182.505 106.590 ;
        RECT 217.360 104.875 217.690 104.890 ;
        RECT 226.560 104.875 226.890 104.890 ;
        RECT 229.780 104.875 230.110 104.890 ;
        RECT 217.360 104.575 230.110 104.875 ;
        RECT 217.360 104.560 217.690 104.575 ;
        RECT 226.560 104.560 226.890 104.575 ;
        RECT 229.780 104.560 230.110 104.575 ;
        RECT 177.625 103.540 179.205 103.870 ;
        RECT 208.620 102.155 208.950 102.170 ;
        RECT 212.760 102.155 213.090 102.170 ;
        RECT 232.540 102.155 232.870 102.170 ;
        RECT 254.160 102.155 254.490 102.170 ;
        RECT 208.620 101.855 254.490 102.155 ;
        RECT 208.620 101.840 208.950 101.855 ;
        RECT 212.760 101.840 213.090 101.855 ;
        RECT 232.540 101.840 232.870 101.855 ;
        RECT 254.160 101.840 254.490 101.855 ;
        RECT 257.840 102.155 258.170 102.170 ;
        RECT 280.840 102.155 281.170 102.170 ;
        RECT 257.840 101.855 281.170 102.155 ;
        RECT 257.840 101.840 258.170 101.855 ;
        RECT 280.840 101.840 281.170 101.855 ;
        RECT 314.335 101.625 314.635 152.405 ;
        RECT 217.360 101.475 217.690 101.490 ;
        RECT 229.780 101.475 230.110 101.490 ;
        RECT 217.360 101.175 230.110 101.475 ;
        RECT 217.360 101.160 217.690 101.175 ;
        RECT 229.780 101.160 230.110 101.175 ;
        RECT 308.900 101.475 309.230 101.490 ;
        RECT 312.335 101.475 314.635 101.625 ;
        RECT 308.900 101.175 314.635 101.475 ;
        RECT 308.900 101.160 309.230 101.175 ;
        RECT 180.925 100.820 182.505 101.150 ;
        RECT 312.335 101.025 314.635 101.175 ;
        RECT 199.880 100.795 200.210 100.810 ;
        RECT 215.060 100.795 215.390 100.810 ;
        RECT 220.580 100.795 220.910 100.810 ;
        RECT 199.880 100.495 220.910 100.795 ;
        RECT 199.880 100.480 200.210 100.495 ;
        RECT 215.060 100.480 215.390 100.495 ;
        RECT 220.580 100.480 220.910 100.495 ;
        RECT 269.340 100.795 269.670 100.810 ;
        RECT 299.240 100.795 299.570 100.810 ;
        RECT 269.340 100.495 299.570 100.795 ;
        RECT 269.340 100.480 269.670 100.495 ;
        RECT 299.240 100.480 299.570 100.495 ;
        RECT 194.360 99.435 194.690 99.450 ;
        RECT 229.320 99.435 229.650 99.450 ;
        RECT 194.360 99.135 229.650 99.435 ;
        RECT 194.360 99.120 194.690 99.135 ;
        RECT 229.320 99.120 229.650 99.135 ;
        RECT 227.940 98.755 228.270 98.770 ;
        RECT 257.380 98.755 257.710 98.770 ;
        RECT 227.940 98.455 257.710 98.755 ;
        RECT 227.940 98.440 228.270 98.455 ;
        RECT 257.380 98.440 257.710 98.455 ;
        RECT 177.625 98.100 179.205 98.430 ;
        RECT 194.820 98.075 195.150 98.090 ;
        RECT 221.500 98.075 221.830 98.090 ;
        RECT 194.820 97.775 221.830 98.075 ;
        RECT 194.820 97.760 195.150 97.775 ;
        RECT 221.500 97.760 221.830 97.775 ;
        RECT 248.180 98.075 248.510 98.090 ;
        RECT 279.920 98.075 280.250 98.090 ;
        RECT 248.180 97.775 280.250 98.075 ;
        RECT 248.180 97.760 248.510 97.775 ;
        RECT 279.920 97.760 280.250 97.775 ;
        RECT 176.880 97.395 177.210 97.410 ;
        RECT 227.940 97.395 228.270 97.410 ;
        RECT 176.880 97.095 228.270 97.395 ;
        RECT 176.880 97.080 177.210 97.095 ;
        RECT 227.940 97.080 228.270 97.095 ;
        RECT 243.580 97.395 243.910 97.410 ;
        RECT 303.380 97.395 303.710 97.410 ;
        RECT 243.580 97.095 303.710 97.395 ;
        RECT 243.580 97.080 243.910 97.095 ;
        RECT 303.380 97.080 303.710 97.095 ;
        RECT 190.220 96.715 190.550 96.730 ;
        RECT 228.400 96.715 228.730 96.730 ;
        RECT 190.220 96.415 228.730 96.715 ;
        RECT 190.220 96.400 190.550 96.415 ;
        RECT 228.400 96.400 228.730 96.415 ;
        RECT 240.820 96.715 241.150 96.730 ;
        RECT 276.240 96.715 276.570 96.730 ;
        RECT 293.720 96.715 294.050 96.730 ;
        RECT 240.820 96.415 294.050 96.715 ;
        RECT 240.820 96.400 241.150 96.415 ;
        RECT 276.240 96.400 276.570 96.415 ;
        RECT 293.720 96.400 294.050 96.415 ;
        RECT 246.800 96.035 247.130 96.050 ;
        RECT 250.020 96.035 250.350 96.050 ;
        RECT 255.080 96.035 255.410 96.050 ;
        RECT 246.800 95.735 255.410 96.035 ;
        RECT 246.800 95.720 247.130 95.735 ;
        RECT 250.020 95.720 250.350 95.735 ;
        RECT 255.080 95.720 255.410 95.735 ;
        RECT 298.780 96.035 299.110 96.050 ;
        RECT 300.160 96.035 300.490 96.050 ;
        RECT 298.780 95.735 300.490 96.035 ;
        RECT 298.780 95.720 299.110 95.735 ;
        RECT 300.160 95.720 300.490 95.735 ;
        RECT 180.925 95.380 182.505 95.710 ;
        RECT 229.320 95.355 229.650 95.370 ;
        RECT 258.760 95.355 259.090 95.370 ;
        RECT 277.160 95.355 277.490 95.370 ;
        RECT 229.320 95.055 277.490 95.355 ;
        RECT 229.320 95.040 229.650 95.055 ;
        RECT 258.760 95.040 259.090 95.055 ;
        RECT 277.160 95.040 277.490 95.055 ;
        RECT 298.780 95.355 299.110 95.370 ;
        RECT 302.000 95.355 302.330 95.370 ;
        RECT 302.920 95.355 303.250 95.370 ;
        RECT 298.780 95.055 303.250 95.355 ;
        RECT 298.780 95.040 299.110 95.055 ;
        RECT 302.000 95.040 302.330 95.055 ;
        RECT 302.920 95.040 303.250 95.055 ;
        RECT 225.180 94.675 225.510 94.690 ;
        RECT 227.940 94.675 228.270 94.690 ;
        RECT 234.840 94.675 235.170 94.690 ;
        RECT 225.180 94.375 235.170 94.675 ;
        RECT 225.180 94.360 225.510 94.375 ;
        RECT 227.940 94.360 228.270 94.375 ;
        RECT 234.840 94.360 235.170 94.375 ;
        RECT 241.280 94.675 241.610 94.690 ;
        RECT 249.100 94.675 249.430 94.690 ;
        RECT 241.280 94.375 249.430 94.675 ;
        RECT 241.280 94.360 241.610 94.375 ;
        RECT 249.100 94.360 249.430 94.375 ;
        RECT 252.780 94.675 253.110 94.690 ;
        RECT 297.860 94.675 298.190 94.690 ;
        RECT 252.780 94.375 298.190 94.675 ;
        RECT 252.780 94.360 253.110 94.375 ;
        RECT 297.860 94.360 298.190 94.375 ;
        RECT 186.080 93.995 186.410 94.010 ;
        RECT 188.840 93.995 189.170 94.010 ;
        RECT 209.080 93.995 209.410 94.010 ;
        RECT 186.080 93.695 209.410 93.995 ;
        RECT 186.080 93.680 186.410 93.695 ;
        RECT 188.840 93.680 189.170 93.695 ;
        RECT 209.080 93.680 209.410 93.695 ;
        RECT 235.300 93.995 235.630 94.010 ;
        RECT 306.140 93.995 306.470 94.010 ;
        RECT 235.300 93.695 306.470 93.995 ;
        RECT 235.300 93.680 235.630 93.695 ;
        RECT 306.140 93.680 306.470 93.695 ;
        RECT 159.185 93.315 161.335 93.465 ;
        RECT 164.000 93.315 164.330 93.330 ;
        RECT 159.185 93.015 164.330 93.315 ;
        RECT 159.185 92.865 161.335 93.015 ;
        RECT 164.000 93.000 164.330 93.015 ;
        RECT 245.880 93.315 246.210 93.330 ;
        RECT 251.400 93.315 251.730 93.330 ;
        RECT 245.880 93.015 251.730 93.315 ;
        RECT 245.880 93.000 246.210 93.015 ;
        RECT 251.400 93.000 251.730 93.015 ;
        RECT 177.625 92.660 179.205 92.990 ;
        RECT 210.460 91.955 210.790 91.970 ;
        RECT 250.480 91.955 250.810 91.970 ;
        RECT 210.460 91.655 250.810 91.955 ;
        RECT 210.460 91.640 210.790 91.655 ;
        RECT 250.480 91.640 250.810 91.655 ;
        RECT 192.060 91.275 192.390 91.290 ;
        RECT 202.640 91.275 202.970 91.290 ;
        RECT 259.680 91.275 260.010 91.290 ;
        RECT 192.060 90.975 260.010 91.275 ;
        RECT 192.060 90.960 192.390 90.975 ;
        RECT 202.640 90.960 202.970 90.975 ;
        RECT 259.680 90.960 260.010 90.975 ;
        RECT 243.580 90.595 243.910 90.610 ;
        RECT 255.080 90.595 255.410 90.610 ;
        RECT 243.580 90.295 255.410 90.595 ;
        RECT 243.580 90.280 243.910 90.295 ;
        RECT 255.080 90.280 255.410 90.295 ;
        RECT 180.925 89.940 182.505 90.270 ;
        RECT 183.780 89.235 184.110 89.250 ;
        RECT 262.900 89.235 263.230 89.250 ;
        RECT 183.780 88.935 263.230 89.235 ;
        RECT 183.780 88.920 184.110 88.935 ;
        RECT 262.900 88.920 263.230 88.935 ;
        RECT 187.000 88.565 187.330 88.570 ;
        RECT 187.000 88.555 187.585 88.565 ;
        RECT 224.720 88.555 225.050 88.570 ;
        RECT 246.800 88.555 247.130 88.570 ;
        RECT 187.000 88.255 187.785 88.555 ;
        RECT 224.720 88.255 247.130 88.555 ;
        RECT 187.000 88.245 187.585 88.255 ;
        RECT 187.000 88.240 187.330 88.245 ;
        RECT 224.720 88.240 225.050 88.255 ;
        RECT 246.800 88.240 247.130 88.255 ;
        RECT 259.220 88.555 259.550 88.570 ;
        RECT 287.740 88.555 288.070 88.570 ;
        RECT 259.220 88.255 288.070 88.555 ;
        RECT 259.220 88.240 259.550 88.255 ;
        RECT 287.740 88.240 288.070 88.255 ;
        RECT 177.625 87.220 179.205 87.550 ;
        RECT 212.300 87.195 212.630 87.210 ;
        RECT 244.500 87.195 244.830 87.210 ;
        RECT 212.300 86.895 244.830 87.195 ;
        RECT 212.300 86.880 212.630 86.895 ;
        RECT 244.500 86.880 244.830 86.895 ;
        RECT 196.200 86.515 196.530 86.530 ;
        RECT 243.580 86.515 243.910 86.530 ;
        RECT 196.200 86.215 243.910 86.515 ;
        RECT 196.200 86.200 196.530 86.215 ;
        RECT 243.580 86.200 243.910 86.215 ;
        RECT 196.660 85.835 196.990 85.850 ;
        RECT 228.400 85.835 228.730 85.850 ;
        RECT 196.660 85.535 228.730 85.835 ;
        RECT 196.660 85.520 196.990 85.535 ;
        RECT 228.400 85.520 228.730 85.535 ;
        RECT 247.720 85.835 248.050 85.850 ;
        RECT 250.480 85.835 250.810 85.850 ;
        RECT 247.720 85.535 250.810 85.835 ;
        RECT 247.720 85.520 248.050 85.535 ;
        RECT 250.480 85.520 250.810 85.535 ;
        RECT 307.520 85.155 307.850 85.170 ;
        RECT 312.335 85.155 314.335 85.305 ;
        RECT 307.520 85.145 314.335 85.155 ;
        RECT 315.070 85.145 315.370 153.575 ;
        RECT 307.520 84.855 315.370 85.145 ;
        RECT 307.520 84.840 307.850 84.855 ;
        RECT 312.335 84.845 315.370 84.855 ;
        RECT 180.925 84.500 182.505 84.830 ;
        RECT 312.335 84.705 314.335 84.845 ;
        RECT 215.060 83.795 215.390 83.810 ;
        RECT 280.380 83.795 280.710 83.810 ;
        RECT 215.060 83.495 280.710 83.795 ;
        RECT 215.060 83.480 215.390 83.495 ;
        RECT 280.380 83.480 280.710 83.495 ;
        RECT 242.660 83.115 242.990 83.130 ;
        RECT 243.325 83.115 243.705 83.125 ;
        RECT 286.360 83.115 286.690 83.130 ;
        RECT 242.660 82.815 286.690 83.115 ;
        RECT 242.660 82.800 242.990 82.815 ;
        RECT 243.325 82.805 243.705 82.815 ;
        RECT 286.360 82.800 286.690 82.815 ;
        RECT 208.620 82.435 208.950 82.450 ;
        RECT 224.720 82.435 225.050 82.450 ;
        RECT 249.100 82.435 249.430 82.450 ;
        RECT 208.620 82.135 249.430 82.435 ;
        RECT 208.620 82.120 208.950 82.135 ;
        RECT 224.720 82.120 225.050 82.135 ;
        RECT 249.100 82.120 249.430 82.135 ;
        RECT 177.625 81.780 179.205 82.110 ;
        RECT 180.100 81.755 180.430 81.770 ;
        RECT 255.540 81.755 255.870 81.770 ;
        RECT 180.100 81.455 255.870 81.755 ;
        RECT 180.100 81.440 180.430 81.455 ;
        RECT 255.540 81.440 255.870 81.455 ;
        RECT 226.560 81.075 226.890 81.090 ;
        RECT 235.300 81.075 235.630 81.090 ;
        RECT 241.740 81.075 242.070 81.090 ;
        RECT 252.320 81.075 252.650 81.090 ;
        RECT 226.560 80.775 252.650 81.075 ;
        RECT 226.560 80.760 226.890 80.775 ;
        RECT 235.300 80.760 235.630 80.775 ;
        RECT 241.740 80.760 242.070 80.775 ;
        RECT 252.320 80.760 252.650 80.775 ;
        RECT 256.920 81.075 257.250 81.090 ;
        RECT 266.120 81.075 266.450 81.090 ;
        RECT 256.920 80.775 266.450 81.075 ;
        RECT 256.920 80.760 257.250 80.775 ;
        RECT 266.120 80.760 266.450 80.775 ;
        RECT 190.680 80.395 191.010 80.410 ;
        RECT 194.565 80.395 194.945 80.405 ;
        RECT 190.680 80.095 194.945 80.395 ;
        RECT 190.680 80.080 191.010 80.095 ;
        RECT 194.565 80.085 194.945 80.095 ;
        RECT 231.620 80.395 231.950 80.410 ;
        RECT 235.045 80.395 235.425 80.405 ;
        RECT 231.620 80.095 235.425 80.395 ;
        RECT 231.620 80.080 231.950 80.095 ;
        RECT 235.045 80.085 235.425 80.095 ;
        RECT 243.580 80.395 243.910 80.410 ;
        RECT 244.245 80.395 244.625 80.405 ;
        RECT 243.580 80.095 244.625 80.395 ;
        RECT 243.580 80.080 243.910 80.095 ;
        RECT 244.245 80.085 244.625 80.095 ;
        RECT 248.180 80.395 248.510 80.410 ;
        RECT 248.845 80.395 249.225 80.405 ;
        RECT 266.120 80.395 266.450 80.410 ;
        RECT 248.180 80.095 249.225 80.395 ;
        RECT 248.180 80.080 248.510 80.095 ;
        RECT 248.845 80.085 249.225 80.095 ;
        RECT 262.685 80.095 266.450 80.395 ;
        RECT 215.520 79.715 215.850 79.730 ;
        RECT 244.500 79.715 244.830 79.730 ;
        RECT 215.520 79.415 244.830 79.715 ;
        RECT 215.520 79.400 215.850 79.415 ;
        RECT 244.500 79.400 244.830 79.415 ;
        RECT 261.060 79.715 261.390 79.730 ;
        RECT 262.685 79.715 262.985 80.095 ;
        RECT 266.120 80.080 266.450 80.095 ;
        RECT 261.060 79.415 262.985 79.715 ;
        RECT 261.060 79.400 261.390 79.415 ;
        RECT 180.925 79.060 182.505 79.390 ;
        RECT 196.660 78.355 196.990 78.370 ;
        RECT 270.260 78.355 270.590 78.370 ;
        RECT 196.660 78.055 270.590 78.355 ;
        RECT 196.660 78.040 196.990 78.055 ;
        RECT 270.260 78.040 270.590 78.055 ;
        RECT 181.020 77.675 181.350 77.690 ;
        RECT 183.320 77.675 183.650 77.690 ;
        RECT 244.040 77.675 244.370 77.690 ;
        RECT 181.020 77.375 244.370 77.675 ;
        RECT 181.020 77.360 181.350 77.375 ;
        RECT 183.320 77.360 183.650 77.375 ;
        RECT 244.040 77.360 244.370 77.375 ;
        RECT 177.625 76.340 179.205 76.670 ;
        RECT 262.440 76.315 262.770 76.330 ;
        RECT 262.440 76.000 262.985 76.315 ;
        RECT 215.060 74.955 215.390 74.970 ;
        RECT 219.660 74.955 219.990 74.970 ;
        RECT 215.060 74.655 219.990 74.955 ;
        RECT 262.685 74.955 262.985 76.000 ;
        RECT 263.360 74.955 263.690 74.970 ;
        RECT 279.000 74.955 279.330 74.970 ;
        RECT 287.740 74.955 288.070 74.970 ;
        RECT 262.685 74.655 288.070 74.955 ;
        RECT 215.060 74.640 215.390 74.655 ;
        RECT 219.660 74.640 219.990 74.655 ;
        RECT 263.360 74.640 263.690 74.655 ;
        RECT 279.000 74.640 279.330 74.655 ;
        RECT 287.740 74.640 288.070 74.655 ;
        RECT 218.280 74.285 218.610 74.290 ;
        RECT 218.280 74.275 218.865 74.285 ;
        RECT 218.055 73.975 218.865 74.275 ;
        RECT 218.280 73.965 218.865 73.975 ;
        RECT 225.640 74.275 225.970 74.290 ;
        RECT 227.480 74.275 227.810 74.290 ;
        RECT 259.680 74.275 260.010 74.290 ;
        RECT 225.640 73.975 260.010 74.275 ;
        RECT 218.280 73.960 218.610 73.965 ;
        RECT 225.640 73.960 225.970 73.975 ;
        RECT 227.480 73.960 227.810 73.975 ;
        RECT 259.680 73.960 260.010 73.975 ;
        RECT 180.925 73.620 182.505 73.950 ;
        RECT 188.840 72.915 189.170 72.930 ;
        RECT 190.220 72.915 190.550 72.930 ;
        RECT 188.840 72.615 190.550 72.915 ;
        RECT 188.840 72.600 189.170 72.615 ;
        RECT 190.220 72.600 190.550 72.615 ;
        RECT 241.740 72.915 242.070 72.930 ;
        RECT 243.325 72.915 243.705 72.925 ;
        RECT 241.740 72.615 243.705 72.915 ;
        RECT 241.740 72.600 242.070 72.615 ;
        RECT 243.325 72.605 243.705 72.615 ;
        RECT 244.245 72.915 244.625 72.925 ;
        RECT 264.740 72.915 265.070 72.930 ;
        RECT 282.220 72.915 282.550 72.930 ;
        RECT 244.245 72.615 282.550 72.915 ;
        RECT 244.245 72.605 244.625 72.615 ;
        RECT 264.740 72.600 265.070 72.615 ;
        RECT 282.220 72.600 282.550 72.615 ;
        RECT 293.260 72.915 293.590 72.930 ;
        RECT 302.920 72.915 303.250 72.930 ;
        RECT 293.260 72.615 303.250 72.915 ;
        RECT 293.260 72.600 293.590 72.615 ;
        RECT 302.920 72.600 303.250 72.615 ;
        RECT 184.700 72.235 185.030 72.250 ;
        RECT 200.800 72.235 201.130 72.250 ;
        RECT 184.700 71.935 201.130 72.235 ;
        RECT 184.700 71.920 185.030 71.935 ;
        RECT 200.800 71.920 201.130 71.935 ;
        RECT 213.220 72.235 213.550 72.250 ;
        RECT 217.820 72.235 218.150 72.250 ;
        RECT 213.220 71.935 218.150 72.235 ;
        RECT 213.220 71.920 213.550 71.935 ;
        RECT 217.820 71.920 218.150 71.935 ;
        RECT 235.045 72.235 235.425 72.245 ;
        RECT 245.880 72.235 246.210 72.250 ;
        RECT 235.045 71.935 246.210 72.235 ;
        RECT 235.045 71.925 235.425 71.935 ;
        RECT 245.880 71.920 246.210 71.935 ;
        RECT 258.300 72.235 258.630 72.250 ;
        RECT 265.660 72.235 265.990 72.250 ;
        RECT 258.300 71.935 265.990 72.235 ;
        RECT 258.300 71.920 258.630 71.935 ;
        RECT 265.660 71.920 265.990 71.935 ;
        RECT 290.960 72.235 291.290 72.250 ;
        RECT 303.380 72.235 303.710 72.250 ;
        RECT 290.960 71.935 303.710 72.235 ;
        RECT 290.960 71.920 291.290 71.935 ;
        RECT 303.380 71.920 303.710 71.935 ;
        RECT 211.380 71.555 211.710 71.570 ;
        RECT 243.120 71.555 243.450 71.570 ;
        RECT 211.380 71.255 243.450 71.555 ;
        RECT 211.380 71.240 211.710 71.255 ;
        RECT 243.120 71.240 243.450 71.255 ;
        RECT 260.140 71.555 260.470 71.570 ;
        RECT 262.900 71.555 263.230 71.570 ;
        RECT 260.140 71.255 263.230 71.555 ;
        RECT 260.140 71.240 260.470 71.255 ;
        RECT 262.900 71.240 263.230 71.255 ;
        RECT 177.625 70.900 179.205 71.230 ;
        RECT 240.820 70.875 241.150 70.890 ;
        RECT 248.180 70.875 248.510 70.890 ;
        RECT 253.240 70.875 253.570 70.890 ;
        RECT 240.820 70.575 253.570 70.875 ;
        RECT 240.820 70.560 241.150 70.575 ;
        RECT 248.180 70.560 248.510 70.575 ;
        RECT 253.240 70.560 253.570 70.575 ;
        RECT 177.800 70.195 178.130 70.210 ;
        RECT 190.220 70.195 190.550 70.210 ;
        RECT 177.800 69.895 190.550 70.195 ;
        RECT 177.800 69.880 178.130 69.895 ;
        RECT 190.220 69.880 190.550 69.895 ;
        RECT 210.920 70.195 211.250 70.210 ;
        RECT 234.840 70.195 235.170 70.210 ;
        RECT 210.920 69.895 235.170 70.195 ;
        RECT 210.920 69.880 211.250 69.895 ;
        RECT 234.840 69.880 235.170 69.895 ;
        RECT 243.580 70.195 243.910 70.210 ;
        RECT 247.260 70.195 247.590 70.210 ;
        RECT 248.640 70.205 248.970 70.210 ;
        RECT 248.640 70.195 249.225 70.205 ;
        RECT 290.040 70.195 290.370 70.210 ;
        RECT 293.260 70.195 293.590 70.210 ;
        RECT 243.580 69.895 247.590 70.195 ;
        RECT 248.435 69.895 293.590 70.195 ;
        RECT 243.580 69.880 243.910 69.895 ;
        RECT 247.260 69.880 247.590 69.895 ;
        RECT 248.640 69.885 249.225 69.895 ;
        RECT 248.640 69.880 248.970 69.885 ;
        RECT 290.040 69.880 290.370 69.895 ;
        RECT 293.260 69.880 293.590 69.895 ;
        RECT 183.780 69.515 184.110 69.530 ;
        RECT 186.080 69.515 186.410 69.530 ;
        RECT 183.780 69.215 186.410 69.515 ;
        RECT 183.780 69.200 184.110 69.215 ;
        RECT 186.080 69.200 186.410 69.215 ;
        RECT 190.680 69.515 191.010 69.530 ;
        RECT 229.780 69.515 230.110 69.530 ;
        RECT 190.680 69.215 230.110 69.515 ;
        RECT 190.680 69.200 191.010 69.215 ;
        RECT 229.780 69.200 230.110 69.215 ;
        RECT 246.340 69.515 246.670 69.530 ;
        RECT 247.005 69.515 247.385 69.525 ;
        RECT 246.340 69.215 247.385 69.515 ;
        RECT 246.340 69.200 246.670 69.215 ;
        RECT 247.005 69.205 247.385 69.215 ;
        RECT 264.280 69.515 264.610 69.530 ;
        RECT 282.680 69.515 283.010 69.530 ;
        RECT 264.280 69.215 283.010 69.515 ;
        RECT 264.280 69.200 264.610 69.215 ;
        RECT 282.680 69.200 283.010 69.215 ;
        RECT 193.900 68.835 194.230 68.850 ;
        RECT 196.200 68.835 196.530 68.850 ;
        RECT 218.280 68.835 218.610 68.850 ;
        RECT 193.900 68.535 218.610 68.835 ;
        RECT 193.900 68.520 194.230 68.535 ;
        RECT 196.200 68.520 196.530 68.535 ;
        RECT 218.280 68.520 218.610 68.535 ;
        RECT 235.300 68.835 235.630 68.850 ;
        RECT 307.980 68.835 308.310 68.850 ;
        RECT 235.300 68.535 308.310 68.835 ;
        RECT 235.300 68.520 235.630 68.535 ;
        RECT 307.980 68.520 308.310 68.535 ;
        RECT 309.360 68.835 309.690 68.850 ;
        RECT 312.335 68.835 314.335 68.985 ;
        RECT 309.360 68.820 314.335 68.835 ;
        RECT 315.845 68.820 316.145 154.625 ;
        RECT 309.360 68.535 316.145 68.820 ;
        RECT 309.360 68.520 309.690 68.535 ;
        RECT 312.335 68.520 316.145 68.535 ;
        RECT 180.925 68.180 182.505 68.510 ;
        RECT 312.335 68.385 314.335 68.520 ;
        RECT 196.660 68.155 196.990 68.170 ;
        RECT 204.480 68.155 204.810 68.170 ;
        RECT 266.580 68.155 266.910 68.170 ;
        RECT 196.660 67.855 266.910 68.155 ;
        RECT 196.660 67.840 196.990 67.855 ;
        RECT 204.480 67.840 204.810 67.855 ;
        RECT 266.580 67.840 266.910 67.855 ;
        RECT 185.620 67.475 185.950 67.490 ;
        RECT 190.680 67.475 191.010 67.490 ;
        RECT 185.620 67.175 191.010 67.475 ;
        RECT 185.620 67.160 185.950 67.175 ;
        RECT 190.680 67.160 191.010 67.175 ;
        RECT 210.000 67.475 210.330 67.490 ;
        RECT 213.680 67.475 214.010 67.490 ;
        RECT 269.340 67.475 269.670 67.490 ;
        RECT 210.000 67.175 269.670 67.475 ;
        RECT 210.000 67.160 210.330 67.175 ;
        RECT 213.680 67.160 214.010 67.175 ;
        RECT 269.340 67.160 269.670 67.175 ;
        RECT 197.120 66.795 197.450 66.810 ;
        RECT 200.800 66.795 201.130 66.810 ;
        RECT 197.120 66.495 201.130 66.795 ;
        RECT 197.120 66.480 197.450 66.495 ;
        RECT 200.800 66.480 201.130 66.495 ;
        RECT 213.680 66.795 214.010 66.810 ;
        RECT 217.360 66.795 217.690 66.810 ;
        RECT 213.680 66.495 217.690 66.795 ;
        RECT 213.680 66.480 214.010 66.495 ;
        RECT 217.360 66.480 217.690 66.495 ;
        RECT 220.580 66.795 220.910 66.810 ;
        RECT 234.840 66.795 235.170 66.810 ;
        RECT 280.380 66.795 280.710 66.810 ;
        RECT 296.020 66.795 296.350 66.810 ;
        RECT 220.580 66.495 222.505 66.795 ;
        RECT 220.580 66.480 220.910 66.495 ;
        RECT 186.080 66.115 186.410 66.130 ;
        RECT 200.340 66.115 200.670 66.130 ;
        RECT 218.280 66.115 218.610 66.130 ;
        RECT 186.080 65.815 218.610 66.115 ;
        RECT 186.080 65.800 186.410 65.815 ;
        RECT 200.340 65.800 200.670 65.815 ;
        RECT 218.280 65.800 218.610 65.815 ;
        RECT 177.625 65.460 179.205 65.790 ;
        RECT 192.520 65.435 192.850 65.450 ;
        RECT 194.360 65.435 194.690 65.450 ;
        RECT 196.660 65.435 196.990 65.450 ;
        RECT 221.500 65.435 221.830 65.450 ;
        RECT 192.520 65.135 221.830 65.435 ;
        RECT 222.205 65.435 222.505 66.495 ;
        RECT 234.840 66.495 296.350 66.795 ;
        RECT 234.840 66.480 235.170 66.495 ;
        RECT 280.380 66.480 280.710 66.495 ;
        RECT 296.020 66.480 296.350 66.495 ;
        RECT 235.760 66.115 236.090 66.130 ;
        RECT 238.980 66.115 239.310 66.130 ;
        RECT 244.500 66.125 244.830 66.130 ;
        RECT 244.245 66.115 244.830 66.125 ;
        RECT 235.760 65.815 239.310 66.115 ;
        RECT 244.045 65.815 244.830 66.115 ;
        RECT 235.760 65.800 236.090 65.815 ;
        RECT 238.980 65.800 239.310 65.815 ;
        RECT 244.245 65.805 244.830 65.815 ;
        RECT 244.500 65.800 244.830 65.805 ;
        RECT 245.880 66.115 246.210 66.130 ;
        RECT 287.740 66.115 288.070 66.130 ;
        RECT 245.880 65.815 288.070 66.115 ;
        RECT 245.880 65.800 246.210 65.815 ;
        RECT 287.740 65.800 288.070 65.815 ;
        RECT 231.160 65.435 231.490 65.450 ;
        RECT 222.205 65.135 231.490 65.435 ;
        RECT 192.520 65.120 192.850 65.135 ;
        RECT 194.360 65.120 194.690 65.135 ;
        RECT 196.660 65.120 196.990 65.135 ;
        RECT 221.500 65.120 221.830 65.135 ;
        RECT 231.160 65.120 231.490 65.135 ;
        RECT 202.180 64.755 202.510 64.770 ;
        RECT 218.280 64.755 218.610 64.770 ;
        RECT 260.600 64.755 260.930 64.770 ;
        RECT 202.180 64.455 217.905 64.755 ;
        RECT 202.180 64.440 202.510 64.455 ;
        RECT 206.780 64.075 207.110 64.090 ;
        RECT 212.760 64.075 213.090 64.090 ;
        RECT 216.900 64.075 217.230 64.090 ;
        RECT 206.780 63.775 217.230 64.075 ;
        RECT 217.605 64.075 217.905 64.455 ;
        RECT 218.280 64.455 260.930 64.755 ;
        RECT 218.280 64.440 218.610 64.455 ;
        RECT 260.600 64.440 260.930 64.455 ;
        RECT 252.320 64.075 252.650 64.090 ;
        RECT 217.605 63.775 252.650 64.075 ;
        RECT 206.780 63.760 207.110 63.775 ;
        RECT 212.760 63.760 213.090 63.775 ;
        RECT 216.900 63.760 217.230 63.775 ;
        RECT 252.320 63.760 252.650 63.775 ;
        RECT 195.740 63.395 196.070 63.410 ;
        RECT 244.040 63.395 244.370 63.410 ;
        RECT 195.740 63.095 244.370 63.395 ;
        RECT 195.740 63.080 196.070 63.095 ;
        RECT 244.040 63.080 244.370 63.095 ;
        RECT 180.925 62.740 182.505 63.070 ;
        RECT 213.220 62.715 213.550 62.730 ;
        RECT 218.740 62.715 219.070 62.730 ;
        RECT 213.220 62.415 219.070 62.715 ;
        RECT 213.220 62.400 213.550 62.415 ;
        RECT 218.740 62.400 219.070 62.415 ;
        RECT 221.500 62.715 221.830 62.730 ;
        RECT 260.140 62.715 260.470 62.730 ;
        RECT 221.500 62.415 260.470 62.715 ;
        RECT 221.500 62.400 221.830 62.415 ;
        RECT 260.140 62.400 260.470 62.415 ;
        RECT 212.300 62.035 212.630 62.050 ;
        RECT 221.960 62.035 222.290 62.050 ;
        RECT 212.300 61.735 222.290 62.035 ;
        RECT 212.300 61.720 212.630 61.735 ;
        RECT 221.960 61.720 222.290 61.735 ;
        RECT 238.980 62.035 239.310 62.050 ;
        RECT 296.480 62.035 296.810 62.050 ;
        RECT 238.980 61.735 296.810 62.035 ;
        RECT 238.980 61.720 239.310 61.735 ;
        RECT 296.480 61.720 296.810 61.735 ;
        RECT 218.485 61.355 218.865 61.365 ;
        RECT 257.380 61.355 257.710 61.370 ;
        RECT 284.520 61.355 284.850 61.370 ;
        RECT 218.485 61.055 284.850 61.355 ;
        RECT 218.485 61.045 218.865 61.055 ;
        RECT 257.380 61.040 257.710 61.055 ;
        RECT 284.520 61.040 284.850 61.055 ;
        RECT 159.335 60.675 161.335 60.825 ;
        RECT 164.000 60.675 164.330 60.690 ;
        RECT 158.335 60.375 164.330 60.675 ;
        RECT 159.335 60.225 161.335 60.375 ;
        RECT 164.000 60.360 164.330 60.375 ;
        RECT 177.625 60.020 179.205 60.350 ;
        RECT 187.205 59.315 187.585 59.325 ;
        RECT 193.900 59.315 194.230 59.330 ;
        RECT 187.205 59.015 194.230 59.315 ;
        RECT 187.205 59.005 187.585 59.015 ;
        RECT 193.900 59.000 194.230 59.015 ;
        RECT 194.565 59.315 194.945 59.325 ;
        RECT 195.280 59.315 195.610 59.330 ;
        RECT 194.565 59.015 195.610 59.315 ;
        RECT 194.565 59.005 194.945 59.015 ;
        RECT 195.280 59.000 195.610 59.015 ;
        RECT 221.500 59.315 221.830 59.330 ;
        RECT 239.900 59.315 240.230 59.330 ;
        RECT 258.300 59.315 258.630 59.330 ;
        RECT 221.500 59.015 258.630 59.315 ;
        RECT 221.500 59.000 221.830 59.015 ;
        RECT 239.900 59.000 240.230 59.015 ;
        RECT 258.300 59.000 258.630 59.015 ;
        RECT 175.960 58.635 176.290 58.650 ;
        RECT 192.520 58.635 192.850 58.650 ;
        RECT 175.960 58.335 192.850 58.635 ;
        RECT 175.960 58.320 176.290 58.335 ;
        RECT 192.520 58.320 192.850 58.335 ;
        RECT 180.925 57.300 182.505 57.630 ;
        RECT 185.620 57.275 185.950 57.290 ;
        RECT 198.040 57.275 198.370 57.290 ;
        RECT 185.620 56.975 198.370 57.275 ;
        RECT 185.620 56.960 185.950 56.975 ;
        RECT 198.040 56.960 198.370 56.975 ;
        RECT 209.540 57.275 209.870 57.290 ;
        RECT 213.680 57.275 214.010 57.290 ;
        RECT 227.480 57.275 227.810 57.290 ;
        RECT 209.540 56.975 227.810 57.275 ;
        RECT 209.540 56.960 209.870 56.975 ;
        RECT 213.680 56.960 214.010 56.975 ;
        RECT 227.480 56.960 227.810 56.975 ;
        RECT 210.460 56.595 210.790 56.610 ;
        RECT 215.980 56.595 216.310 56.610 ;
        RECT 210.460 56.295 216.310 56.595 ;
        RECT 210.460 56.280 210.790 56.295 ;
        RECT 215.980 56.280 216.310 56.295 ;
        RECT 177.625 54.580 179.205 54.910 ;
        RECT 183.780 54.555 184.110 54.570 ;
        RECT 246.800 54.555 247.130 54.570 ;
        RECT 183.780 54.255 247.130 54.555 ;
        RECT 183.780 54.240 184.110 54.255 ;
        RECT 246.800 54.240 247.130 54.255 ;
        RECT 175.960 53.875 176.290 53.890 ;
        RECT 244.500 53.875 244.830 53.890 ;
        RECT 175.960 53.575 244.830 53.875 ;
        RECT 175.960 53.560 176.290 53.575 ;
        RECT 244.500 53.560 244.830 53.575 ;
        RECT 245.880 53.875 246.210 53.890 ;
        RECT 278.540 53.875 278.870 53.890 ;
        RECT 245.880 53.575 278.870 53.875 ;
        RECT 245.880 53.560 246.210 53.575 ;
        RECT 278.540 53.560 278.870 53.575 ;
        RECT 309.360 52.515 309.690 52.530 ;
        RECT 312.335 52.515 314.335 52.665 ;
        RECT 309.360 52.505 314.335 52.515 ;
        RECT 316.545 52.505 316.845 155.650 ;
        RECT 309.360 52.215 316.845 52.505 ;
        RECT 309.360 52.200 309.690 52.215 ;
        RECT 312.335 52.205 316.845 52.215 ;
        RECT 180.925 51.860 182.505 52.190 ;
        RECT 312.335 52.065 314.335 52.205 ;
        RECT 204.020 50.475 204.350 50.490 ;
        RECT 259.220 50.475 259.550 50.490 ;
        RECT 204.020 50.175 259.550 50.475 ;
        RECT 204.020 50.160 204.350 50.175 ;
        RECT 259.220 50.160 259.550 50.175 ;
        RECT 177.625 49.140 179.205 49.470 ;
        RECT 180.925 46.420 182.505 46.750 ;
        RECT 177.625 43.700 179.205 44.030 ;
        RECT 180.925 40.980 182.505 41.310 ;
        RECT 177.625 38.260 179.205 38.590 ;
        RECT 316.555 36.345 316.955 36.545 ;
        RECT 308.900 36.195 309.230 36.210 ;
        RECT 312.335 36.195 316.955 36.345 ;
        RECT 308.900 35.895 316.955 36.195 ;
        RECT 308.900 35.880 309.230 35.895 ;
        RECT 180.925 35.540 182.505 35.870 ;
        RECT 312.335 35.745 316.955 35.895 ;
        RECT 177.625 32.820 179.205 33.150 ;
        RECT 180.925 30.100 182.505 30.430 ;
        RECT 159.335 28.035 161.335 28.185 ;
        RECT 164.000 28.035 164.330 28.050 ;
        RECT 157.560 27.735 164.330 28.035 ;
        RECT 159.335 27.585 161.335 27.735 ;
        RECT 164.000 27.720 164.330 27.735 ;
        RECT 177.625 27.380 179.205 27.710 ;
        RECT 180.925 24.660 182.505 24.990 ;
        RECT 177.625 21.940 179.205 22.270 ;
        RECT 247.005 19.875 247.385 19.885 ;
        RECT 312.335 19.875 314.335 20.025 ;
        RECT 247.005 19.845 314.335 19.875 ;
        RECT 317.375 19.845 317.675 156.780 ;
        RECT 318.485 36.545 318.785 157.875 ;
        RECT 318.085 35.745 318.785 36.545 ;
        RECT 247.005 19.575 317.675 19.845 ;
        RECT 247.005 19.565 247.385 19.575 ;
        RECT 180.925 19.220 182.505 19.550 ;
        RECT 312.335 19.545 317.675 19.575 ;
        RECT 312.335 19.425 314.335 19.545 ;
        RECT 177.625 16.500 179.205 16.830 ;
        RECT 180.925 13.780 182.505 14.110 ;
      LAYER met4 ;
        RECT 23.260 224.760 23.310 225.560 ;
        RECT 23.610 224.760 23.660 225.560 ;
        RECT 45.340 224.760 45.390 225.560 ;
        RECT 45.690 224.760 45.740 225.560 ;
        RECT 65.010 225.310 65.510 225.710 ;
        RECT 125.730 225.360 126.530 225.760 ;
        RECT 59.490 224.760 59.990 225.160 ;
        RECT 67.770 224.760 68.270 225.110 ;
        RECT 129.395 225.050 130.195 225.100 ;
        RECT 75.700 224.760 75.750 224.860 ;
        RECT 76.050 224.760 76.100 224.860 ;
        RECT 78.810 224.760 78.945 224.860 ;
        RECT 15.030 224.460 15.330 224.760 ;
        RECT 17.790 224.460 18.090 224.760 ;
        RECT 20.550 224.460 20.850 224.760 ;
        RECT 26.070 224.460 26.370 224.760 ;
        RECT 28.830 224.460 29.130 224.760 ;
        RECT 31.590 224.460 31.890 224.760 ;
        RECT 34.350 224.460 34.650 224.760 ;
        RECT 37.110 224.460 37.410 224.760 ;
        RECT 39.870 224.460 40.170 224.760 ;
        RECT 42.630 224.460 42.930 224.760 ;
        RECT 48.150 224.460 48.450 224.760 ;
        RECT 50.910 224.460 51.210 224.760 ;
        RECT 53.670 224.460 53.970 224.760 ;
        RECT 56.430 224.460 56.730 224.760 ;
        RECT 3.600 224.060 56.730 224.460 ;
        RECT 61.950 224.560 62.250 224.760 ;
        RECT 67.470 224.710 68.270 224.760 ;
        RECT 61.950 224.160 62.750 224.560 ;
        RECT 70.230 224.510 70.530 224.760 ;
        RECT 70.230 224.110 71.030 224.510 ;
        RECT 1.000 220.760 1.800 221.560 ;
        RECT 3.600 220.760 5.200 224.060 ;
        RECT 72.990 223.910 73.290 224.760 ;
        RECT 75.700 224.060 76.100 224.760 ;
        RECT 78.510 224.060 78.945 224.760 ;
        RECT 83.980 224.760 84.030 224.860 ;
        RECT 84.330 224.760 84.380 224.860 ;
        RECT 83.980 224.060 84.380 224.760 ;
        RECT 86.740 224.760 86.790 224.860 ;
        RECT 87.090 224.760 87.140 224.860 ;
        RECT 86.740 224.060 87.140 224.760 ;
        RECT 92.260 224.760 92.310 224.860 ;
        RECT 92.610 224.760 92.660 224.860 ;
        RECT 128.490 224.760 130.195 225.050 ;
        RECT 92.260 224.060 92.660 224.760 ;
        RECT 95.070 224.450 95.370 224.760 ;
        RECT 97.830 224.450 98.130 224.760 ;
        RECT 100.590 224.450 100.890 224.760 ;
        RECT 103.350 224.450 103.650 224.760 ;
        RECT 106.110 224.450 106.410 224.760 ;
        RECT 108.870 224.615 109.170 224.760 ;
        RECT 72.990 223.510 73.790 223.910 ;
        RECT 95.020 223.650 95.420 224.450 ;
        RECT 97.780 223.650 98.180 224.450 ;
        RECT 100.540 223.650 100.940 224.450 ;
        RECT 103.300 223.650 103.700 224.450 ;
        RECT 106.060 223.650 106.460 224.450 ;
        RECT 108.865 224.215 109.665 224.615 ;
        RECT 6.200 221.180 109.540 222.780 ;
        RECT 111.630 221.515 111.930 224.760 ;
        RECT 114.390 222.115 114.690 224.760 ;
        RECT 117.150 222.715 117.450 224.760 ;
        RECT 119.910 223.315 120.210 224.760 ;
        RECT 122.670 223.915 122.970 224.760 ;
        RECT 128.190 224.750 130.195 224.760 ;
        RECT 129.395 224.700 130.195 224.750 ;
        RECT 122.670 223.615 149.190 223.915 ;
        RECT 119.910 223.015 145.160 223.315 ;
        RECT 117.150 222.415 141.130 222.715 ;
        RECT 114.390 221.815 137.100 222.115 ;
        RECT 136.800 221.515 137.100 221.815 ;
        RECT 140.830 221.515 141.130 222.415 ;
        RECT 144.860 221.515 145.160 223.015 ;
        RECT 148.890 221.515 149.190 223.615 ;
      LAYER met4 ;
        RECT 255.465 221.585 317.065 223.185 ;
      LAYER met4 ;
        RECT 111.630 221.215 133.120 221.515 ;
        RECT 6.200 220.760 7.800 221.180 ;
        RECT 10.550 218.590 105.040 220.190 ;
        RECT 7.800 211.890 11.170 215.090 ;
        RECT 43.720 211.890 45.320 215.090 ;
        RECT 103.440 211.240 105.040 218.590 ;
        RECT 106.340 219.305 109.540 221.180 ;
        RECT 132.720 220.715 133.120 221.215 ;
        RECT 136.750 220.715 137.150 221.515 ;
        RECT 140.780 220.715 141.180 221.515 ;
        RECT 144.810 220.715 145.210 221.515 ;
        RECT 148.840 220.715 149.240 221.515 ;
        RECT 106.340 217.705 151.230 219.305 ;
        RECT 106.340 217.515 109.540 217.705 ;
        RECT 106.415 211.240 108.015 213.740 ;
        RECT 150.830 211.240 248.550 212.040 ;
        RECT 27.080 209.940 53.660 210.740 ;
        RECT 27.080 209.640 27.570 209.940 ;
        RECT 16.115 199.365 25.725 208.975 ;
        RECT 16.115 196.975 16.715 199.365 ;
        RECT 16.115 187.365 25.725 196.975 ;
        RECT 16.115 184.975 16.715 187.365 ;
        RECT 16.115 175.365 25.725 184.975 ;
        RECT 16.115 172.975 16.715 175.365 ;
        RECT 16.115 163.365 25.725 172.975 ;
        RECT 16.115 160.975 16.715 163.365 ;
        RECT 16.115 151.365 25.725 160.975 ;
        RECT 16.115 150.210 16.715 151.365 ;
        RECT 27.080 150.970 27.565 209.640 ;
        RECT 28.915 199.365 38.525 208.975 ;
        RECT 37.925 196.975 38.525 199.365 ;
        RECT 28.915 187.365 38.525 196.975 ;
        RECT 52.860 188.465 53.660 209.940 ;
        RECT 103.440 209.640 248.550 211.240 ;
        RECT 150.830 208.840 248.550 209.640 ;
        RECT 173.605 199.585 175.205 208.840 ;
        RECT 177.405 189.425 177.735 189.755 ;
        RECT 110.530 187.540 156.765 189.140 ;
        RECT 37.925 184.975 38.525 187.365 ;
        RECT 28.915 175.365 38.525 184.975 ;
        RECT 37.925 172.975 38.525 175.365 ;
        RECT 28.915 163.365 38.525 172.975 ;
        RECT 51.950 184.940 103.750 186.540 ;
        RECT 51.950 169.890 53.550 184.940 ;
        RECT 57.020 177.390 109.070 178.990 ;
        RECT 153.565 178.210 156.765 187.540 ;
        RECT 175.565 183.985 175.895 184.315 ;
        RECT 175.580 179.555 175.880 183.985 ;
        RECT 177.420 179.555 177.720 189.425 ;
        RECT 179.245 186.025 179.575 186.355 ;
        RECT 175.565 179.225 175.895 179.555 ;
        RECT 177.405 179.225 177.735 179.555 ;
        RECT 179.260 178.875 179.560 186.025 ;
        RECT 179.245 178.545 179.575 178.875 ;
        RECT 151.155 175.010 156.765 178.210 ;
        RECT 180.670 176.770 182.270 201.730 ;
        RECT 182.925 183.985 183.255 184.315 ;
        RECT 182.940 180.235 183.240 183.985 ;
        RECT 182.925 179.905 183.255 180.235 ;
        RECT 183.970 178.360 185.570 201.730 ;
        RECT 192.115 199.585 193.715 208.840 ;
        RECT 210.625 199.585 212.225 208.840 ;
        RECT 229.135 199.585 230.735 208.840 ;
        RECT 190.285 185.345 190.615 185.675 ;
        RECT 182.860 176.770 185.570 178.360 ;
        RECT 190.300 177.515 190.600 185.345 ;
        RECT 212.365 184.665 212.695 184.995 ;
        RECT 212.380 179.555 212.680 184.665 ;
        RECT 212.365 179.225 212.695 179.555 ;
        RECT 190.285 177.185 190.615 177.515 ;
        RECT 51.950 168.290 58.420 169.890 ;
        RECT 37.925 160.975 38.525 163.365 ;
        RECT 28.915 151.365 38.525 160.975 ;
        RECT 153.565 168.200 156.765 175.010 ;
        RECT 182.860 168.200 184.460 176.770 ;
        RECT 201.370 168.200 202.970 178.360 ;
        RECT 219.880 168.200 221.480 178.360 ;
        RECT 238.390 168.200 239.990 178.360 ;
        RECT 153.565 165.000 240.760 168.200 ;
        RECT 111.685 158.165 112.085 158.565 ;
        RECT 105.385 157.765 112.085 158.165 ;
        RECT 105.385 157.365 105.785 157.765 ;
        RECT 109.415 156.565 109.815 156.965 ;
        RECT 113.085 156.565 113.485 156.965 ;
        RECT 109.415 156.165 113.485 156.565 ;
        RECT 37.925 150.210 38.525 151.365 ;
        RECT 16.115 149.410 46.630 150.210 ;
        RECT 51.575 145.090 73.495 148.290 ;
        RECT 9.490 135.030 17.100 142.640 ;
        RECT 18.455 142.175 20.750 142.975 ;
        RECT 13.385 130.025 14.185 135.030 ;
        RECT 18.455 134.695 18.935 142.175 ;
        RECT 20.350 141.375 20.750 142.175 ;
        RECT 61.980 135.495 62.780 135.895 ;
        RECT 61.980 135.095 140.370 135.495 ;
        RECT 22.615 133.320 80.925 134.120 ;
        RECT 20.650 131.810 21.050 132.210 ;
        RECT 137.945 131.810 138.345 132.210 ;
        RECT 20.650 131.410 138.345 131.810 ;
        RECT 139.120 130.025 139.520 132.990 ;
        RECT 13.385 129.625 139.520 130.025 ;
        RECT 16.805 128.710 139.520 129.110 ;
        RECT 65.865 124.285 67.465 127.485 ;
        RECT 121.565 124.285 123.165 127.485 ;
        RECT 139.120 125.690 139.520 128.710 ;
        RECT 139.970 125.690 140.370 135.095 ;
        RECT 140.940 131.390 142.100 132.990 ;
        RECT 140.940 125.060 141.340 131.390 ;
        RECT 131.145 124.660 141.340 125.060 ;
        RECT 103.315 121.565 118.965 123.165 ;
        RECT 109.865 107.965 118.715 109.565 ;
        RECT 63.315 103.465 74.365 105.065 ;
        RECT 105.965 103.615 118.565 105.215 ;
        RECT 131.145 98.015 131.545 124.660 ;
        RECT 153.565 124.090 156.765 165.000 ;
        RECT 142.760 122.490 156.765 124.090 ;
        RECT 153.565 114.150 156.765 122.490 ;
        RECT 139.355 113.350 156.765 114.150 ;
        RECT 245.350 113.705 248.550 208.840 ;
      LAYER met4 ;
        RECT 255.465 207.185 257.065 221.585 ;
      LAYER met4 ;
        RECT 257.065 219.185 271.465 221.585 ;
      LAYER met4 ;
        RECT 271.465 219.585 277.065 221.585 ;
      LAYER met4 ;
        RECT 277.065 219.585 279.465 221.585 ;
      LAYER met4 ;
        RECT 279.465 219.585 285.065 221.585 ;
      LAYER met4 ;
        RECT 285.065 219.585 289.465 221.585 ;
      LAYER met4 ;
        RECT 289.465 219.585 293.065 221.585 ;
      LAYER met4 ;
        RECT 293.065 219.585 297.465 221.585 ;
      LAYER met4 ;
        RECT 297.465 219.585 301.065 221.585 ;
      LAYER met4 ;
        RECT 257.065 209.585 259.465 219.185 ;
      LAYER met4 ;
        RECT 259.465 217.585 269.065 219.185 ;
        RECT 259.465 211.185 261.065 217.585 ;
      LAYER met4 ;
        RECT 261.065 211.185 267.465 217.585 ;
      LAYER met4 ;
        RECT 267.465 211.185 269.065 217.585 ;
        RECT 259.465 209.585 269.065 211.185 ;
      LAYER met4 ;
        RECT 269.065 209.585 271.465 219.185 ;
      LAYER met4 ;
        RECT 271.465 215.185 273.065 219.585 ;
      LAYER met4 ;
        RECT 273.065 217.185 279.465 219.585 ;
      LAYER met4 ;
        RECT 279.465 217.185 283.065 219.585 ;
      LAYER met4 ;
        RECT 283.065 217.185 289.465 219.585 ;
      LAYER met4 ;
        RECT 289.465 217.185 291.065 219.585 ;
      LAYER met4 ;
        RECT 291.065 219.185 299.465 219.585 ;
        RECT 291.065 217.585 295.465 219.185 ;
      LAYER met4 ;
        RECT 295.465 217.585 297.065 219.185 ;
      LAYER met4 ;
        RECT 297.065 217.585 299.465 219.185 ;
        RECT 291.065 217.185 299.465 217.585 ;
        RECT 273.065 215.585 275.465 217.185 ;
      LAYER met4 ;
        RECT 275.465 215.585 291.065 217.185 ;
      LAYER met4 ;
        RECT 291.065 215.585 293.465 217.185 ;
      LAYER met4 ;
        RECT 293.465 215.585 295.065 217.185 ;
      LAYER met4 ;
        RECT 295.065 215.585 299.465 217.185 ;
        RECT 273.065 215.185 277.465 215.585 ;
      LAYER met4 ;
        RECT 271.465 213.585 275.065 215.185 ;
      LAYER met4 ;
        RECT 275.065 213.585 277.465 215.185 ;
      LAYER met4 ;
        RECT 277.465 213.585 281.065 215.585 ;
      LAYER met4 ;
        RECT 281.065 213.585 285.465 215.585 ;
      LAYER met4 ;
        RECT 285.465 213.585 287.065 215.585 ;
      LAYER met4 ;
        RECT 287.065 213.585 289.465 215.585 ;
      LAYER met4 ;
        RECT 289.465 215.185 291.065 215.585 ;
      LAYER met4 ;
        RECT 291.065 215.185 299.465 215.585 ;
      LAYER met4 ;
        RECT 289.465 213.585 293.065 215.185 ;
      LAYER met4 ;
        RECT 293.065 213.585 299.465 215.185 ;
        RECT 257.065 207.185 271.465 209.585 ;
      LAYER met4 ;
        RECT 271.465 207.185 273.065 213.585 ;
      LAYER met4 ;
        RECT 273.065 211.185 279.465 213.585 ;
      LAYER met4 ;
        RECT 255.465 205.585 273.065 207.185 ;
      LAYER met4 ;
        RECT 273.065 205.585 275.465 211.185 ;
      LAYER met4 ;
        RECT 255.465 199.185 257.065 205.585 ;
      LAYER met4 ;
        RECT 257.065 201.585 261.465 205.585 ;
      LAYER met4 ;
        RECT 261.465 203.185 263.065 205.585 ;
      LAYER met4 ;
        RECT 263.065 203.185 265.465 205.585 ;
      LAYER met4 ;
        RECT 265.465 203.585 269.065 205.585 ;
      LAYER met4 ;
        RECT 269.065 205.185 275.465 205.585 ;
      LAYER met4 ;
        RECT 275.465 205.185 277.065 211.185 ;
      LAYER met4 ;
        RECT 277.065 207.585 279.465 211.185 ;
      LAYER met4 ;
        RECT 279.465 207.585 281.065 213.585 ;
      LAYER met4 ;
        RECT 281.065 213.185 299.465 213.585 ;
      LAYER met4 ;
        RECT 299.465 213.185 301.065 219.585 ;
      LAYER met4 ;
        RECT 301.065 219.185 315.465 221.585 ;
        RECT 281.065 207.585 283.465 213.185 ;
      LAYER met4 ;
        RECT 283.465 211.185 285.065 213.185 ;
      LAYER met4 ;
        RECT 285.065 211.585 295.465 213.185 ;
      LAYER met4 ;
        RECT 295.465 211.585 301.065 213.185 ;
      LAYER met4 ;
        RECT 285.065 211.185 297.465 211.585 ;
      LAYER met4 ;
        RECT 283.465 209.585 287.065 211.185 ;
      LAYER met4 ;
        RECT 287.065 209.585 289.465 211.185 ;
      LAYER met4 ;
        RECT 289.465 209.585 295.065 211.185 ;
      LAYER met4 ;
        RECT 295.065 209.585 297.465 211.185 ;
      LAYER met4 ;
        RECT 297.465 209.585 301.065 211.585 ;
      LAYER met4 ;
        RECT 301.065 209.585 303.465 219.185 ;
      LAYER met4 ;
        RECT 303.465 217.585 313.065 219.185 ;
        RECT 303.465 211.185 305.065 217.585 ;
      LAYER met4 ;
        RECT 305.065 211.185 311.465 217.585 ;
      LAYER met4 ;
        RECT 311.465 211.185 313.065 217.585 ;
        RECT 303.465 209.585 313.065 211.185 ;
      LAYER met4 ;
        RECT 313.065 209.585 315.465 219.185 ;
      LAYER met4 ;
        RECT 283.465 207.585 285.065 209.585 ;
      LAYER met4 ;
        RECT 285.065 209.185 291.465 209.585 ;
        RECT 285.065 207.585 287.465 209.185 ;
        RECT 277.065 207.185 287.465 207.585 ;
      LAYER met4 ;
        RECT 287.465 207.185 289.065 209.185 ;
      LAYER met4 ;
        RECT 289.065 207.585 291.465 209.185 ;
      LAYER met4 ;
        RECT 291.465 207.585 293.065 209.585 ;
      LAYER met4 ;
        RECT 293.065 209.185 299.465 209.585 ;
        RECT 293.065 207.585 295.465 209.185 ;
        RECT 277.065 205.585 281.465 207.185 ;
      LAYER met4 ;
        RECT 281.465 205.585 283.065 207.185 ;
      LAYER met4 ;
        RECT 283.065 205.585 285.465 207.185 ;
      LAYER met4 ;
        RECT 285.465 205.585 289.065 207.185 ;
      LAYER met4 ;
        RECT 289.065 205.585 295.465 207.585 ;
      LAYER met4 ;
        RECT 295.465 205.585 297.065 209.185 ;
      LAYER met4 ;
        RECT 297.065 205.585 299.465 209.185 ;
      LAYER met4 ;
        RECT 299.465 207.185 301.065 209.585 ;
      LAYER met4 ;
        RECT 301.065 207.185 315.465 209.585 ;
      LAYER met4 ;
        RECT 315.465 207.185 317.065 221.585 ;
        RECT 299.465 205.585 317.065 207.185 ;
      LAYER met4 ;
        RECT 277.065 205.185 287.465 205.585 ;
      LAYER met4 ;
        RECT 287.465 205.185 289.065 205.585 ;
      LAYER met4 ;
        RECT 289.065 205.185 299.465 205.585 ;
      LAYER met4 ;
        RECT 299.465 205.185 301.065 205.585 ;
      LAYER met4 ;
        RECT 269.065 203.585 273.465 205.185 ;
      LAYER met4 ;
        RECT 273.465 203.585 279.065 205.185 ;
      LAYER met4 ;
        RECT 279.065 203.585 283.465 205.185 ;
      LAYER met4 ;
        RECT 283.465 203.585 285.065 205.185 ;
      LAYER met4 ;
        RECT 285.065 203.585 287.465 205.185 ;
      LAYER met4 ;
        RECT 287.465 203.585 295.065 205.185 ;
      LAYER met4 ;
        RECT 295.065 203.585 297.465 205.185 ;
      LAYER met4 ;
        RECT 297.465 203.585 301.065 205.185 ;
      LAYER met4 ;
        RECT 301.065 203.585 307.465 205.585 ;
      LAYER met4 ;
        RECT 307.465 203.585 309.065 205.585 ;
      LAYER met4 ;
        RECT 309.065 203.585 313.465 205.585 ;
      LAYER met4 ;
        RECT 313.465 203.585 317.065 205.585 ;
        RECT 265.465 203.185 267.065 203.585 ;
      LAYER met4 ;
        RECT 267.065 203.185 277.465 203.585 ;
      LAYER met4 ;
        RECT 261.465 201.585 267.065 203.185 ;
      LAYER met4 ;
        RECT 267.065 201.585 269.465 203.185 ;
      LAYER met4 ;
        RECT 269.465 201.585 271.065 203.185 ;
      LAYER met4 ;
        RECT 271.065 201.585 277.465 203.185 ;
        RECT 257.065 201.185 277.465 201.585 ;
      LAYER met4 ;
        RECT 277.465 201.185 279.065 203.585 ;
      LAYER met4 ;
        RECT 279.065 203.185 287.465 203.585 ;
      LAYER met4 ;
        RECT 287.465 203.185 289.065 203.585 ;
      LAYER met4 ;
        RECT 289.065 203.185 297.465 203.585 ;
      LAYER met4 ;
        RECT 297.465 203.185 299.065 203.585 ;
      LAYER met4 ;
        RECT 299.065 203.185 315.465 203.585 ;
        RECT 279.065 201.585 285.465 203.185 ;
      LAYER met4 ;
        RECT 285.465 201.585 289.065 203.185 ;
      LAYER met4 ;
        RECT 289.065 201.585 295.465 203.185 ;
      LAYER met4 ;
        RECT 295.465 201.585 299.065 203.185 ;
      LAYER met4 ;
        RECT 299.065 201.585 303.465 203.185 ;
      LAYER met4 ;
        RECT 303.465 201.585 307.065 203.185 ;
      LAYER met4 ;
        RECT 257.065 199.185 271.465 201.185 ;
      LAYER met4 ;
        RECT 271.465 199.185 273.065 201.185 ;
      LAYER met4 ;
        RECT 273.065 199.585 275.465 201.185 ;
      LAYER met4 ;
        RECT 275.465 199.585 279.065 201.185 ;
      LAYER met4 ;
        RECT 279.065 199.585 287.465 201.585 ;
      LAYER met4 ;
        RECT 287.465 201.185 289.065 201.585 ;
      LAYER met4 ;
        RECT 289.065 201.185 305.465 201.585 ;
      LAYER met4 ;
        RECT 287.465 199.585 291.065 201.185 ;
      LAYER met4 ;
        RECT 291.065 199.585 299.465 201.185 ;
      LAYER met4 ;
        RECT 299.465 199.585 301.065 201.185 ;
      LAYER met4 ;
        RECT 301.065 199.585 305.465 201.185 ;
        RECT 273.065 199.185 287.465 199.585 ;
      LAYER met4 ;
        RECT 287.465 199.185 289.065 199.585 ;
      LAYER met4 ;
        RECT 289.065 199.185 305.465 199.585 ;
      LAYER met4 ;
        RECT 305.465 199.185 307.065 201.585 ;
      LAYER met4 ;
        RECT 307.065 201.185 315.465 203.185 ;
      LAYER met4 ;
        RECT 315.465 201.185 317.065 203.585 ;
      LAYER met4 ;
        RECT 307.065 199.185 313.465 201.185 ;
      LAYER met4 ;
        RECT 255.465 195.185 259.065 199.185 ;
      LAYER met4 ;
        RECT 259.065 197.585 261.465 199.185 ;
        POLYGON 261.465 199.185 261.770 199.185 261.465 198.880 ;
      LAYER met4 ;
        RECT 261.770 198.880 273.065 199.185 ;
        RECT 261.465 197.585 273.065 198.880 ;
      LAYER met4 ;
        RECT 273.065 197.585 285.465 199.185 ;
      LAYER met4 ;
        RECT 285.465 197.585 289.065 199.185 ;
      LAYER met4 ;
        RECT 289.065 197.585 291.465 199.185 ;
      LAYER met4 ;
        RECT 291.465 197.585 293.065 199.185 ;
      LAYER met4 ;
        RECT 293.065 197.585 301.465 199.185 ;
      LAYER met4 ;
        RECT 301.465 197.585 309.065 199.185 ;
      LAYER met4 ;
        RECT 309.065 197.585 313.465 199.185 ;
      LAYER met4 ;
        RECT 313.465 197.585 317.065 201.185 ;
      LAYER met4 ;
        RECT 259.065 195.585 265.465 197.585 ;
      LAYER met4 ;
        RECT 265.465 195.585 267.065 197.585 ;
      LAYER met4 ;
        RECT 267.065 197.185 287.465 197.585 ;
      LAYER met4 ;
        RECT 287.465 197.185 289.065 197.585 ;
      LAYER met4 ;
        RECT 289.065 197.185 303.465 197.585 ;
        RECT 267.065 195.585 275.465 197.185 ;
        RECT 259.065 195.185 275.465 195.585 ;
      LAYER met4 ;
        RECT 275.465 195.185 277.065 197.185 ;
      LAYER met4 ;
        RECT 277.065 195.185 281.465 197.185 ;
      LAYER met4 ;
        RECT 281.465 195.585 285.065 197.185 ;
      LAYER met4 ;
        RECT 285.065 195.585 287.465 197.185 ;
      LAYER met4 ;
        RECT 255.465 193.585 263.065 195.185 ;
      LAYER met4 ;
        RECT 263.065 193.585 269.465 195.185 ;
      LAYER met4 ;
        RECT 269.465 193.585 273.065 195.185 ;
      LAYER met4 ;
        RECT 273.065 193.585 275.465 195.185 ;
      LAYER met4 ;
        RECT 255.465 191.585 259.065 193.585 ;
      LAYER met4 ;
        RECT 259.065 193.185 275.465 193.585 ;
        RECT 259.065 191.585 263.465 193.185 ;
      LAYER met4 ;
        RECT 263.465 191.585 269.065 193.185 ;
      LAYER met4 ;
        RECT 269.065 191.585 275.465 193.185 ;
      LAYER met4 ;
        RECT 255.465 189.185 257.065 191.585 ;
      LAYER met4 ;
        RECT 257.065 191.185 263.465 191.585 ;
        RECT 257.065 189.585 259.465 191.185 ;
      LAYER met4 ;
        RECT 259.465 189.585 261.065 191.185 ;
      LAYER met4 ;
        RECT 261.065 189.585 263.465 191.185 ;
      LAYER met4 ;
        RECT 263.465 189.585 267.065 191.585 ;
      LAYER met4 ;
        RECT 267.065 191.185 275.465 191.585 ;
      LAYER met4 ;
        RECT 275.465 191.185 279.065 195.185 ;
      LAYER met4 ;
        RECT 267.065 189.585 269.465 191.185 ;
      LAYER met4 ;
        RECT 269.465 189.585 271.065 191.185 ;
      LAYER met4 ;
        RECT 271.065 189.585 273.465 191.185 ;
      LAYER met4 ;
        RECT 273.465 189.585 279.065 191.185 ;
      LAYER met4 ;
        RECT 279.065 189.585 281.465 195.185 ;
      LAYER met4 ;
        RECT 281.465 191.185 283.065 195.585 ;
      LAYER met4 ;
        RECT 283.065 191.585 287.465 195.585 ;
      LAYER met4 ;
        RECT 287.465 191.585 291.065 197.185 ;
      LAYER met4 ;
        RECT 291.065 191.585 293.465 197.185 ;
      LAYER met4 ;
        RECT 293.465 193.185 295.065 197.185 ;
      LAYER met4 ;
        RECT 295.065 195.185 303.465 197.185 ;
      LAYER met4 ;
        RECT 303.465 195.185 307.065 197.585 ;
      LAYER met4 ;
        RECT 307.065 197.185 315.465 197.585 ;
        RECT 295.065 193.185 299.465 195.185 ;
      LAYER met4 ;
        RECT 299.465 193.585 307.065 195.185 ;
        RECT 299.465 193.185 301.065 193.585 ;
        RECT 293.465 191.585 301.065 193.185 ;
      LAYER met4 ;
        RECT 301.065 191.585 303.465 193.585 ;
      LAYER met4 ;
        RECT 303.465 191.585 307.065 193.585 ;
      LAYER met4 ;
        RECT 307.065 191.585 309.465 197.185 ;
      LAYER met4 ;
        RECT 309.465 195.185 311.065 197.185 ;
      LAYER met4 ;
        RECT 311.065 195.185 315.465 197.185 ;
      LAYER met4 ;
        RECT 315.465 195.185 317.065 197.585 ;
        RECT 309.465 193.585 317.065 195.185 ;
      LAYER met4 ;
        RECT 283.065 191.185 297.465 191.585 ;
      LAYER met4 ;
        RECT 281.465 189.585 287.065 191.185 ;
      LAYER met4 ;
        RECT 257.065 189.185 263.465 189.585 ;
      LAYER met4 ;
        RECT 263.465 189.185 265.065 189.585 ;
      LAYER met4 ;
        RECT 265.065 189.185 273.465 189.585 ;
      LAYER met4 ;
        RECT 255.465 185.585 259.065 189.185 ;
      LAYER met4 ;
        RECT 259.065 185.585 261.465 189.185 ;
      LAYER met4 ;
        RECT 261.465 187.890 265.065 189.185 ;
        RECT 261.465 187.585 264.760 187.890 ;
        POLYGON 264.760 187.890 265.065 187.890 264.760 187.585 ;
      LAYER met4 ;
        RECT 265.065 187.585 267.465 189.185 ;
      LAYER met4 ;
        RECT 267.465 187.585 269.065 189.185 ;
      LAYER met4 ;
        RECT 269.065 187.585 273.465 189.185 ;
      LAYER met4 ;
        RECT 261.465 185.585 263.065 187.585 ;
      LAYER met4 ;
        RECT 263.065 187.185 273.465 187.585 ;
      LAYER met4 ;
        RECT 273.465 187.185 275.065 189.585 ;
      LAYER met4 ;
        RECT 275.065 187.585 277.465 189.585 ;
      LAYER met4 ;
        RECT 277.465 189.185 279.065 189.585 ;
      LAYER met4 ;
        RECT 279.065 189.185 285.465 189.585 ;
      LAYER met4 ;
        RECT 277.465 187.585 281.065 189.185 ;
      LAYER met4 ;
        RECT 281.065 187.585 285.465 189.185 ;
      LAYER met4 ;
        RECT 285.465 187.585 287.065 189.585 ;
      LAYER met4 ;
        RECT 287.065 189.185 297.465 191.185 ;
        RECT 287.065 187.585 289.465 189.185 ;
        RECT 263.065 185.585 269.465 187.185 ;
      LAYER met4 ;
        RECT 269.465 185.585 275.065 187.185 ;
      LAYER met4 ;
        RECT 275.065 185.585 279.465 187.585 ;
      LAYER met4 ;
        RECT 279.465 185.585 281.065 187.585 ;
      LAYER met4 ;
        RECT 281.065 187.185 289.465 187.585 ;
      LAYER met4 ;
        RECT 289.465 187.185 291.065 189.185 ;
      LAYER met4 ;
        RECT 291.065 187.585 293.465 189.185 ;
      LAYER met4 ;
        RECT 293.465 187.585 295.065 189.185 ;
      LAYER met4 ;
        RECT 295.065 187.585 297.465 189.185 ;
        RECT 291.065 187.185 297.465 187.585 ;
      LAYER met4 ;
        RECT 297.465 187.185 299.065 191.585 ;
      LAYER met4 ;
        RECT 299.065 189.185 303.465 191.585 ;
      LAYER met4 ;
        RECT 303.465 189.185 305.065 191.585 ;
      LAYER met4 ;
        RECT 305.065 191.185 309.465 191.585 ;
      LAYER met4 ;
        RECT 309.465 191.185 311.065 193.585 ;
      LAYER met4 ;
        RECT 311.065 191.185 315.465 193.585 ;
      LAYER met4 ;
        RECT 315.465 191.185 317.065 193.585 ;
      LAYER met4 ;
        RECT 305.065 189.585 307.465 191.185 ;
      LAYER met4 ;
        RECT 307.465 189.585 317.065 191.185 ;
      LAYER met4 ;
        RECT 305.065 189.185 309.465 189.585 ;
        RECT 299.065 187.585 301.465 189.185 ;
      LAYER met4 ;
        RECT 301.465 187.585 307.065 189.185 ;
      LAYER met4 ;
        RECT 307.065 187.585 309.465 189.185 ;
      LAYER met4 ;
        RECT 309.465 187.585 313.065 189.585 ;
      LAYER met4 ;
        RECT 313.065 187.585 315.465 189.585 ;
        RECT 281.065 185.585 287.465 187.185 ;
      LAYER met4 ;
        RECT 287.465 185.585 293.065 187.185 ;
      LAYER met4 ;
        RECT 293.065 185.585 295.465 187.185 ;
      LAYER met4 ;
        RECT 255.465 183.185 257.065 185.585 ;
      LAYER met4 ;
        RECT 257.065 185.185 273.465 185.585 ;
      LAYER met4 ;
        RECT 273.465 185.185 275.065 185.585 ;
      LAYER met4 ;
        RECT 275.065 185.185 287.465 185.585 ;
        RECT 257.065 183.185 259.465 185.185 ;
      LAYER met4 ;
        RECT 259.465 183.185 261.065 185.185 ;
      LAYER met4 ;
        RECT 261.065 183.185 263.465 185.185 ;
      LAYER met4 ;
        RECT 263.465 183.185 265.065 185.185 ;
      LAYER met4 ;
        RECT 265.065 183.185 273.465 185.185 ;
      LAYER met4 ;
        RECT 273.465 183.585 277.065 185.185 ;
      LAYER met4 ;
        RECT 277.065 183.585 283.465 185.185 ;
      LAYER met4 ;
        RECT 255.465 181.585 265.065 183.185 ;
      LAYER met4 ;
        RECT 265.065 181.585 267.465 183.185 ;
      LAYER met4 ;
        RECT 267.465 181.585 271.065 183.185 ;
      LAYER met4 ;
        RECT 271.065 181.585 273.465 183.185 ;
      LAYER met4 ;
        RECT 255.465 179.185 257.065 181.585 ;
      LAYER met4 ;
        RECT 257.065 179.185 259.465 181.585 ;
      LAYER met4 ;
        RECT 259.465 179.185 265.065 181.585 ;
      LAYER met4 ;
        RECT 265.065 181.185 273.465 181.585 ;
      LAYER met4 ;
        RECT 273.465 181.185 275.065 183.585 ;
      LAYER met4 ;
        RECT 275.065 183.185 283.465 183.585 ;
        RECT 275.065 181.185 279.465 183.185 ;
      LAYER met4 ;
        RECT 279.465 181.185 281.065 183.185 ;
      LAYER met4 ;
        RECT 281.065 181.185 283.465 183.185 ;
      LAYER met4 ;
        RECT 283.465 181.185 285.065 185.185 ;
      LAYER met4 ;
        RECT 285.065 183.585 287.465 185.185 ;
      LAYER met4 ;
        RECT 287.465 183.585 289.065 185.585 ;
      LAYER met4 ;
        RECT 289.065 183.585 295.465 185.585 ;
      LAYER met4 ;
        RECT 295.465 185.185 299.065 187.185 ;
      LAYER met4 ;
        RECT 299.065 185.585 303.465 187.585 ;
      LAYER met4 ;
        RECT 303.465 185.585 307.065 187.585 ;
      LAYER met4 ;
        RECT 307.065 185.585 315.465 187.585 ;
        RECT 299.065 185.185 315.465 185.585 ;
      LAYER met4 ;
        RECT 295.465 183.585 303.065 185.185 ;
      LAYER met4 ;
        RECT 303.065 183.585 307.465 185.185 ;
        RECT 285.065 183.185 299.465 183.585 ;
        RECT 285.065 181.585 293.465 183.185 ;
      LAYER met4 ;
        RECT 293.465 181.585 295.065 183.185 ;
      LAYER met4 ;
        RECT 295.065 181.585 299.465 183.185 ;
      LAYER met4 ;
        RECT 299.465 181.585 301.065 183.585 ;
      LAYER met4 ;
        RECT 301.065 183.185 307.465 183.585 ;
      LAYER met4 ;
        RECT 307.465 183.185 311.065 185.185 ;
      LAYER met4 ;
        RECT 311.065 183.185 315.465 185.185 ;
      LAYER met4 ;
        RECT 315.465 183.185 317.065 189.585 ;
      LAYER met4 ;
        RECT 301.065 181.585 303.465 183.185 ;
      LAYER met4 ;
        RECT 303.465 181.585 305.065 183.185 ;
      LAYER met4 ;
        RECT 305.065 181.585 307.465 183.185 ;
      LAYER met4 ;
        RECT 307.465 181.585 317.065 183.185 ;
      LAYER met4 ;
        RECT 285.065 181.185 307.465 181.585 ;
        RECT 265.065 179.185 271.465 181.185 ;
      LAYER met4 ;
        RECT 271.465 179.585 275.065 181.185 ;
      LAYER met4 ;
        RECT 275.065 179.585 277.465 181.185 ;
      LAYER met4 ;
        RECT 277.465 179.890 293.065 181.185 ;
      LAYER met4 ;
        POLYGON 277.465 179.890 277.770 179.585 277.465 179.585 ;
      LAYER met4 ;
        RECT 277.770 179.585 293.065 179.890 ;
        RECT 271.465 179.185 273.065 179.585 ;
        RECT 255.465 177.585 273.065 179.185 ;
        RECT 255.465 163.185 257.065 177.585 ;
      LAYER met4 ;
        RECT 257.065 175.185 271.465 177.585 ;
      LAYER met4 ;
        RECT 271.465 175.185 273.065 177.585 ;
      LAYER met4 ;
        RECT 273.065 177.185 281.465 179.585 ;
      LAYER met4 ;
        RECT 281.465 177.185 285.065 179.585 ;
      LAYER met4 ;
        RECT 285.065 177.185 287.465 179.585 ;
      LAYER met4 ;
        RECT 287.465 179.185 293.065 179.585 ;
      LAYER met4 ;
        RECT 293.065 179.185 307.465 181.185 ;
      LAYER met4 ;
        RECT 287.465 177.585 295.065 179.185 ;
        RECT 287.465 177.185 289.065 177.585 ;
      LAYER met4 ;
        RECT 273.065 175.585 277.465 177.185 ;
      LAYER met4 ;
        RECT 277.465 175.585 289.065 177.185 ;
      LAYER met4 ;
        RECT 289.065 175.585 293.465 177.585 ;
      LAYER met4 ;
        RECT 293.465 177.185 295.065 177.585 ;
      LAYER met4 ;
        RECT 295.065 177.185 299.465 179.185 ;
      LAYER met4 ;
        RECT 299.465 177.585 305.065 179.185 ;
      LAYER met4 ;
        RECT 305.065 177.585 307.465 179.185 ;
      LAYER met4 ;
        RECT 307.465 177.585 309.065 181.585 ;
      LAYER met4 ;
        RECT 309.065 177.585 315.465 181.585 ;
      LAYER met4 ;
        RECT 293.465 175.585 297.065 177.185 ;
      LAYER met4 ;
        RECT 273.065 175.185 279.465 175.585 ;
        RECT 257.065 165.585 259.465 175.185 ;
      LAYER met4 ;
        RECT 259.465 173.585 269.065 175.185 ;
        RECT 259.465 167.185 261.065 173.585 ;
      LAYER met4 ;
        RECT 261.065 167.185 267.465 173.585 ;
      LAYER met4 ;
        RECT 267.465 167.185 269.065 173.585 ;
        RECT 259.465 165.585 269.065 167.185 ;
      LAYER met4 ;
        RECT 269.065 165.585 271.465 175.185 ;
      LAYER met4 ;
        RECT 271.465 173.585 277.065 175.185 ;
      LAYER met4 ;
        RECT 277.065 173.585 279.465 175.185 ;
      LAYER met4 ;
        RECT 279.465 173.585 285.065 175.585 ;
      LAYER met4 ;
        RECT 285.065 175.185 295.465 175.585 ;
      LAYER met4 ;
        RECT 271.465 171.585 275.065 173.585 ;
      LAYER met4 ;
        RECT 275.065 173.185 279.465 173.585 ;
      LAYER met4 ;
        RECT 279.465 173.185 281.065 173.585 ;
      LAYER met4 ;
        RECT 275.065 171.585 277.465 173.185 ;
      LAYER met4 ;
        RECT 277.465 171.585 281.065 173.185 ;
      LAYER met4 ;
        RECT 281.065 171.585 283.465 173.585 ;
      LAYER met4 ;
        RECT 283.465 173.185 285.065 173.585 ;
      LAYER met4 ;
        RECT 285.065 173.185 289.465 175.185 ;
      LAYER met4 ;
        RECT 289.465 173.585 293.065 175.185 ;
      LAYER met4 ;
        RECT 293.065 173.585 295.465 175.185 ;
      LAYER met4 ;
        RECT 289.465 173.185 291.065 173.585 ;
      LAYER met4 ;
        RECT 291.065 173.185 295.465 173.585 ;
      LAYER met4 ;
        RECT 295.465 173.185 297.065 175.585 ;
      LAYER met4 ;
        RECT 297.065 173.585 299.465 177.185 ;
      LAYER met4 ;
        RECT 299.465 175.185 301.065 177.585 ;
      LAYER met4 ;
        RECT 301.065 175.185 303.465 177.585 ;
      LAYER met4 ;
        RECT 303.465 175.185 305.065 177.585 ;
      LAYER met4 ;
        RECT 305.065 177.185 315.465 177.585 ;
      LAYER met4 ;
        RECT 315.465 177.185 317.065 181.585 ;
      LAYER met4 ;
        RECT 305.065 175.585 309.465 177.185 ;
      LAYER met4 ;
        RECT 309.465 175.585 311.065 177.185 ;
      LAYER met4 ;
        RECT 311.065 175.585 313.465 177.185 ;
        RECT 305.065 175.185 313.465 175.585 ;
      LAYER met4 ;
        RECT 313.465 175.185 317.065 177.185 ;
        RECT 299.465 173.585 305.065 175.185 ;
      LAYER met4 ;
        RECT 305.065 173.585 307.465 175.185 ;
      LAYER met4 ;
        RECT 283.465 171.585 291.065 173.185 ;
      LAYER met4 ;
        RECT 291.065 171.585 293.465 173.185 ;
      LAYER met4 ;
        RECT 293.465 171.890 297.065 173.185 ;
      LAYER met4 ;
        POLYGON 293.465 171.890 293.770 171.585 293.465 171.585 ;
      LAYER met4 ;
        RECT 293.770 171.585 297.065 171.890 ;
        RECT 271.465 169.185 273.065 171.585 ;
      LAYER met4 ;
        RECT 273.065 171.185 283.465 171.585 ;
        RECT 273.065 169.585 275.465 171.185 ;
      LAYER met4 ;
        RECT 275.465 169.585 277.065 171.185 ;
      LAYER met4 ;
        RECT 277.065 169.585 283.465 171.185 ;
        RECT 273.065 169.185 283.465 169.585 ;
      LAYER met4 ;
        RECT 271.465 167.585 275.065 169.185 ;
      LAYER met4 ;
        RECT 275.065 167.585 279.465 169.185 ;
        RECT 257.065 163.185 271.465 165.585 ;
      LAYER met4 ;
        RECT 271.465 163.185 273.065 167.585 ;
      LAYER met4 ;
        RECT 273.065 167.185 279.465 167.585 ;
      LAYER met4 ;
        RECT 279.465 167.185 281.065 169.185 ;
      LAYER met4 ;
        RECT 281.065 167.585 283.465 169.185 ;
      LAYER met4 ;
        RECT 283.465 167.585 289.065 171.585 ;
      LAYER met4 ;
        RECT 289.065 169.585 295.465 171.585 ;
      LAYER met4 ;
        RECT 295.465 171.185 297.065 171.585 ;
      LAYER met4 ;
        RECT 297.065 171.185 307.465 173.585 ;
      LAYER met4 ;
        RECT 307.465 173.185 309.065 175.185 ;
      LAYER met4 ;
        RECT 309.065 173.585 311.465 175.185 ;
      LAYER met4 ;
        RECT 311.465 173.585 317.065 175.185 ;
      LAYER met4 ;
        RECT 309.065 173.185 315.465 173.585 ;
      LAYER met4 ;
        RECT 295.465 169.585 301.065 171.185 ;
      LAYER met4 ;
        RECT 301.065 169.585 307.465 171.185 ;
      LAYER met4 ;
        RECT 307.465 169.585 311.065 173.185 ;
      LAYER met4 ;
        RECT 311.065 171.185 315.465 173.185 ;
      LAYER met4 ;
        RECT 315.465 171.185 317.065 173.585 ;
      LAYER met4 ;
        RECT 311.065 169.585 313.465 171.185 ;
      LAYER met4 ;
        RECT 313.465 169.585 317.065 171.185 ;
      LAYER met4 ;
        RECT 289.065 169.185 297.465 169.585 ;
        RECT 289.065 167.585 293.465 169.185 ;
        RECT 273.065 165.585 275.465 167.185 ;
      LAYER met4 ;
        RECT 275.465 165.585 281.065 167.185 ;
      LAYER met4 ;
        RECT 281.065 165.585 293.465 167.585 ;
      LAYER met4 ;
        RECT 293.465 167.185 295.065 169.185 ;
      LAYER met4 ;
        RECT 295.065 167.585 297.465 169.185 ;
      LAYER met4 ;
        RECT 297.465 167.585 299.065 169.585 ;
      LAYER met4 ;
        RECT 299.065 169.185 315.465 169.585 ;
        RECT 299.065 167.585 301.465 169.185 ;
        RECT 295.065 167.185 301.465 167.585 ;
        RECT 273.065 163.185 277.465 165.585 ;
      LAYER met4 ;
        RECT 277.465 163.185 279.065 165.585 ;
      LAYER met4 ;
        RECT 279.065 165.185 293.465 165.585 ;
        RECT 279.065 163.185 281.465 165.185 ;
      LAYER met4 ;
        RECT 281.465 163.185 283.065 165.185 ;
      LAYER met4 ;
        RECT 283.065 163.185 287.465 165.185 ;
      LAYER met4 ;
        RECT 287.465 163.185 289.065 165.185 ;
      LAYER met4 ;
        RECT 289.065 163.185 293.465 165.185 ;
      LAYER met4 ;
        RECT 293.465 163.185 297.065 167.185 ;
      LAYER met4 ;
        RECT 297.065 165.585 301.465 167.185 ;
      LAYER met4 ;
        RECT 301.465 165.585 305.065 169.185 ;
      LAYER met4 ;
        RECT 305.065 167.585 311.465 169.185 ;
      LAYER met4 ;
        RECT 311.465 167.585 313.065 169.185 ;
      LAYER met4 ;
        RECT 313.065 167.585 315.465 169.185 ;
        RECT 305.065 167.185 315.465 167.585 ;
      LAYER met4 ;
        RECT 315.465 167.185 317.065 169.585 ;
      LAYER met4 ;
        RECT 305.065 165.585 307.465 167.185 ;
      LAYER met4 ;
        RECT 307.465 165.585 311.065 167.185 ;
      LAYER met4 ;
        RECT 297.065 165.185 309.465 165.585 ;
        RECT 297.065 163.185 305.465 165.185 ;
      LAYER met4 ;
        RECT 305.465 163.185 307.065 165.185 ;
      LAYER met4 ;
        RECT 307.065 163.185 309.465 165.185 ;
      LAYER met4 ;
        RECT 309.465 163.185 311.065 165.585 ;
      LAYER met4 ;
        RECT 311.065 163.185 313.465 167.185 ;
      LAYER met4 ;
        RECT 313.465 163.185 317.065 167.185 ;
        RECT 255.465 161.585 317.065 163.185 ;
      LAYER met4 ;
        RECT 100.115 96.415 132.145 98.015 ;
        RECT 97.165 93.265 124.815 94.865 ;
        RECT 43.135 78.605 52.745 82.655 ;
        RECT 56.135 78.605 65.745 82.655 ;
        RECT 69.135 78.605 78.745 82.655 ;
        RECT 82.135 78.605 91.745 82.655 ;
        RECT 95.135 78.605 104.745 82.655 ;
        RECT 130.545 78.605 132.145 96.415 ;
        RECT 38.470 77.005 132.145 78.605 ;
        RECT 38.470 63.590 39.745 77.005 ;
        RECT 43.135 73.045 52.745 77.005 ;
        RECT 56.135 73.045 65.745 77.005 ;
        RECT 69.135 73.045 78.745 77.005 ;
        RECT 82.135 73.045 91.745 77.005 ;
        RECT 95.135 73.045 104.745 77.005 ;
        RECT 42.800 71.180 108.800 71.690 ;
        RECT 133.525 71.180 135.125 110.315 ;
        RECT 42.800 69.580 135.125 71.180 ;
        RECT 42.800 69.190 108.800 69.580 ;
        RECT 43.135 63.590 52.745 67.835 ;
        RECT 56.135 63.590 65.745 67.835 ;
        RECT 69.135 63.590 78.745 67.835 ;
        RECT 82.135 63.590 91.745 67.835 ;
        RECT 95.135 63.590 104.745 67.835 ;
        RECT 38.470 61.990 104.745 63.590 ;
        RECT 43.135 58.225 52.745 61.990 ;
        RECT 56.135 58.225 65.745 61.990 ;
        RECT 69.135 58.225 78.745 61.990 ;
        RECT 82.135 58.225 91.745 61.990 ;
        RECT 95.135 58.225 104.745 61.990 ;
        RECT 12.915 45.565 92.315 47.165 ;
        RECT 65.765 42.615 117.715 44.215 ;
        RECT 68.865 40.015 120.815 41.615 ;
        RECT 72.095 9.265 82.535 10.865 ;
        RECT 153.565 8.890 156.765 113.350 ;
        RECT 179.925 110.505 293.305 113.705 ;
        RECT 179.925 106.665 181.525 110.505 ;
        RECT 177.615 13.705 179.215 106.665 ;
        RECT 179.925 103.110 182.515 106.665 ;
        RECT 217.185 103.110 218.785 110.505 ;
        RECT 254.445 103.110 256.045 110.505 ;
        RECT 291.705 103.110 293.305 110.505 ;
        RECT 180.915 13.705 182.515 103.110 ;
        RECT 187.230 88.240 187.560 88.570 ;
        RECT 187.245 59.330 187.545 88.240 ;
        RECT 243.350 82.800 243.680 83.130 ;
        RECT 194.590 80.080 194.920 80.410 ;
        RECT 235.070 80.080 235.400 80.410 ;
        RECT 194.605 59.330 194.905 80.080 ;
        RECT 218.510 73.960 218.840 74.290 ;
        RECT 218.525 61.370 218.825 73.960 ;
        RECT 235.085 72.250 235.385 80.080 ;
        RECT 243.365 72.930 243.665 82.800 ;
        RECT 244.270 80.080 244.600 80.410 ;
        RECT 248.870 80.080 249.200 80.410 ;
        RECT 244.285 72.930 244.585 80.080 ;
        RECT 243.350 72.600 243.680 72.930 ;
        RECT 244.270 72.600 244.600 72.930 ;
        RECT 235.070 71.920 235.400 72.250 ;
        RECT 244.285 66.130 244.585 72.600 ;
        RECT 248.885 70.210 249.185 80.080 ;
        RECT 248.870 69.880 249.200 70.210 ;
        RECT 247.030 69.200 247.360 69.530 ;
        RECT 244.270 65.800 244.600 66.130 ;
        RECT 218.510 61.040 218.840 61.370 ;
        RECT 187.230 59.000 187.560 59.330 ;
        RECT 194.590 59.000 194.920 59.330 ;
        RECT 247.045 19.890 247.345 69.200 ;
        RECT 247.030 19.560 247.360 19.890 ;
        RECT 198.555 8.890 200.155 16.285 ;
        RECT 235.815 8.890 237.415 16.285 ;
        RECT 273.075 8.890 274.675 16.285 ;
        RECT 310.335 8.890 311.935 16.285 ;
        RECT 14.965 5.690 16.565 8.890 ;
        RECT 128.160 5.690 311.935 8.890 ;
        RECT 97.530 1.000 98.430 2.125 ;
        RECT 116.850 1.750 132.465 2.650 ;
        RECT 136.170 1.750 152.360 2.650 ;
        RECT 116.850 1.000 117.750 1.750 ;
        RECT 136.170 1.000 137.070 1.750 ;
  END
END tt_um_cw_vref
END LIBRARY

